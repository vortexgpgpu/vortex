module VX_tex_format #(
    parameter CORE_ID = 0
) (
    // TODO
)   
    `UNUSED_PARAM (CORE_ID)
    
    // TODO

endmodule