`include "VX_platform.vh"

`TRACING_OFF
module VX_mem_streamer #(
    parameter NUM_REQS = 1
    // TODO
) (
    input  wire clk,
    input  wire reset
    // TODO
  );

    // TODO
    
endmodule
`TRACING_ON