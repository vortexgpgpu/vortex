# Copyright (c) 1993 - 2019 ARM Limited. All Rights Reserved.
# Use of this Software is subject to the terms and conditions of the
# applicable license agreement with ARM Limited.

# PhyVGen V 8.8.0
# ARM Version r0p0
# Creation Date: Sun Oct 13 11:08:55 2019


# Memory Configuration:
# ~~~~~~~~~~~~~~~~~~~~~
#  -activity_factor 50 -atf off -back_biasing off -bits 128 -bmux on
# -bus_notation on -check_instname on -diodes on -drive 6 -ema on -frequency
# 1.0 -instname rf2_32x128_wm1 -left_bus_delim "[" -mux 2 -mvt LL -name_case
# upper -pipeline off -power_gating off -power_type otc -pwr_gnd_rename
# vddpe:VDDPE,vddce:VDDCE,vsse:VSSE -rcols 2 -redundancy off -retention on
# -right_bus_delim "]" -rrows 0 -ser none -site_def off -top_layer m5-m10
# -words 32 -wp_size 1 -write_mask on -write_thru off -corners
# ff_0p99v_0p99v_m40c,ss_0p81v_0p81v_125c,tt_0p81v_0p81v_0c
# 

VERSION 5.8 ;
BUSBITCHARS "[]" ;
MACRO rf2_32x128_wm1
	FOREIGN rf2_32x128_wm1 0 0 ;
	SYMMETRY X Y ;
	SIZE 21.975 BY 414.86 ;
	CLASS BLOCK ;
	PIN AA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 191.27 0.25 191.37 ;
			LAYER	M2 ;
			RECT	0 191.27 0.25 191.37 ;
			LAYER	M3 ;
			RECT	0 191.27 0.25 191.37 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[0]

	PIN AA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 194.3 0.25 194.4 ;
			LAYER	M2 ;
			RECT	0 194.3 0.25 194.4 ;
			LAYER	M3 ;
			RECT	0 194.3 0.25 194.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[1]

	PIN AA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 197.33 0.25 197.43 ;
			LAYER	M2 ;
			RECT	0 197.33 0.25 197.43 ;
			LAYER	M3 ;
			RECT	0 197.33 0.25 197.43 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[2]

	PIN AA[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 198.875 0.25 198.975 ;
			LAYER	M2 ;
			RECT	0 198.875 0.25 198.975 ;
			LAYER	M3 ;
			RECT	0 198.875 0.25 198.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[3]

	PIN AA[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 201.905 0.25 202.005 ;
			LAYER	M2 ;
			RECT	0 201.905 0.25 202.005 ;
			LAYER	M3 ;
			RECT	0 201.905 0.25 202.005 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[4]

	PIN AB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 224.185 0.25 224.285 ;
			LAYER	M2 ;
			RECT	0 224.185 0.25 224.285 ;
			LAYER	M3 ;
			RECT	0 224.185 0.25 224.285 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[0]

	PIN AB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 220.96 0.25 221.06 ;
			LAYER	M2 ;
			RECT	0 220.96 0.25 221.06 ;
			LAYER	M3 ;
			RECT	0 220.96 0.25 221.06 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[1]

	PIN AB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 218.125 0.25 218.225 ;
			LAYER	M2 ;
			RECT	0 218.125 0.25 218.225 ;
			LAYER	M3 ;
			RECT	0 218.125 0.25 218.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[2]

	PIN AB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 216.58 0.25 216.68 ;
			LAYER	M2 ;
			RECT	0 216.58 0.25 216.68 ;
			LAYER	M3 ;
			RECT	0 216.58 0.25 216.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[3]

	PIN AB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 213.55 0.25 213.65 ;
			LAYER	M2 ;
			RECT	0 213.55 0.25 213.65 ;
			LAYER	M3 ;
			RECT	0 213.55 0.25 213.65 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[4]

	PIN AYA[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 191.675 0.25 191.775 ;
			LAYER	M2 ;
			RECT	0 191.675 0.25 191.775 ;
			LAYER	M3 ;
			RECT	0 191.675 0.25 191.775 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[0]

	PIN AYA[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 194.705 0.25 194.805 ;
			LAYER	M2 ;
			RECT	0 194.705 0.25 194.805 ;
			LAYER	M3 ;
			RECT	0 194.705 0.25 194.805 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[1]

	PIN AYA[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 197.735 0.25 197.835 ;
			LAYER	M2 ;
			RECT	0 197.735 0.25 197.835 ;
			LAYER	M3 ;
			RECT	0 197.735 0.25 197.835 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[2]

	PIN AYA[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 198.5 0.25 198.6 ;
			LAYER	M2 ;
			RECT	0 198.5 0.25 198.6 ;
			LAYER	M3 ;
			RECT	0 198.5 0.25 198.6 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[3]

	PIN AYA[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 201.705 0.25 201.805 ;
			LAYER	M2 ;
			RECT	0 201.705 0.25 201.805 ;
			LAYER	M3 ;
			RECT	0 201.705 0.25 201.805 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[4]

	PIN AYB[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 223.78 0.25 223.88 ;
			LAYER	M2 ;
			RECT	0 223.78 0.25 223.88 ;
			LAYER	M3 ;
			RECT	0 223.78 0.25 223.88 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[0]

	PIN AYB[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 220.75 0.25 220.85 ;
			LAYER	M2 ;
			RECT	0 220.75 0.25 220.85 ;
			LAYER	M3 ;
			RECT	0 220.75 0.25 220.85 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[1]

	PIN AYB[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 217.75 0.25 217.85 ;
			LAYER	M2 ;
			RECT	0 217.75 0.25 217.85 ;
			LAYER	M3 ;
			RECT	0 217.75 0.25 217.85 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[2]

	PIN AYB[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 216.985 0.25 217.085 ;
			LAYER	M2 ;
			RECT	0 216.985 0.25 217.085 ;
			LAYER	M3 ;
			RECT	0 216.985 0.25 217.085 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[3]

	PIN AYB[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 213.925 0.25 214.025 ;
			LAYER	M2 ;
			RECT	0 213.925 0.25 214.025 ;
			LAYER	M3 ;
			RECT	0 213.925 0.25 214.025 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[4]

	PIN CENA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 188.51 0.25 188.61 ;
			LAYER	M2 ;
			RECT	0 188.51 0.25 188.61 ;
			LAYER	M3 ;
			RECT	0 188.51 0.25 188.61 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENA

	PIN CENB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 228.705 0.25 228.805 ;
			LAYER	M2 ;
			RECT	0 228.705 0.25 228.805 ;
			LAYER	M3 ;
			RECT	0 228.705 0.25 228.805 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENB

	PIN CENYA
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 187.1 0.25 187.2 ;
			LAYER	M2 ;
			RECT	0 187.1 0.25 187.2 ;
			LAYER	M3 ;
			RECT	0 187.1 0.25 187.2 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENYA

	PIN CENYB
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 229.25 0.25 229.35 ;
			LAYER	M2 ;
			RECT	0 229.25 0.25 229.35 ;
			LAYER	M3 ;
			RECT	0 229.25 0.25 229.35 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENYB

	PIN CLKA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 198.13 0.25 198.23 ;
			LAYER	M2 ;
			RECT	0 198.13 0.25 198.23 ;
			LAYER	M3 ;
			RECT	0 198.13 0.25 198.23 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CLKA

	PIN CLKB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 218.78 0.25 218.88 ;
			LAYER	M2 ;
			RECT	0 218.78 0.25 218.88 ;
			LAYER	M3 ;
			RECT	0 218.78 0.25 218.88 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CLKB

	PIN COLLDISN
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 206.3 0.25 206.4 ;
			LAYER	M2 ;
			RECT	0 206.3 0.25 206.4 ;
			LAYER	M3 ;
			RECT	0 206.3 0.25 206.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END COLLDISN

	PIN DB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 2.195 0.25 2.295 ;
			LAYER	M2 ;
			RECT	0 2.195 0.25 2.295 ;
			LAYER	M3 ;
			RECT	0 2.195 0.25 2.295 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[0]

	PIN DB[100]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 334.805 0.25 334.905 ;
			LAYER	M2 ;
			RECT	0 334.805 0.25 334.905 ;
			LAYER	M3 ;
			RECT	0 334.805 0.25 334.905 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[100]

	PIN DB[101]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 337.685 0.25 337.785 ;
			LAYER	M2 ;
			RECT	0 337.685 0.25 337.785 ;
			LAYER	M3 ;
			RECT	0 337.685 0.25 337.785 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[101]

	PIN DB[102]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 340.565 0.25 340.665 ;
			LAYER	M2 ;
			RECT	0 340.565 0.25 340.665 ;
			LAYER	M3 ;
			RECT	0 340.565 0.25 340.665 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[102]

	PIN DB[103]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 343.445 0.25 343.545 ;
			LAYER	M2 ;
			RECT	0 343.445 0.25 343.545 ;
			LAYER	M3 ;
			RECT	0 343.445 0.25 343.545 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[103]

	PIN DB[104]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 346.325 0.25 346.425 ;
			LAYER	M2 ;
			RECT	0 346.325 0.25 346.425 ;
			LAYER	M3 ;
			RECT	0 346.325 0.25 346.425 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[104]

	PIN DB[105]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 349.205 0.25 349.305 ;
			LAYER	M2 ;
			RECT	0 349.205 0.25 349.305 ;
			LAYER	M3 ;
			RECT	0 349.205 0.25 349.305 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[105]

	PIN DB[106]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 352.085 0.25 352.185 ;
			LAYER	M2 ;
			RECT	0 352.085 0.25 352.185 ;
			LAYER	M3 ;
			RECT	0 352.085 0.25 352.185 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[106]

	PIN DB[107]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 354.965 0.25 355.065 ;
			LAYER	M2 ;
			RECT	0 354.965 0.25 355.065 ;
			LAYER	M3 ;
			RECT	0 354.965 0.25 355.065 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[107]

	PIN DB[108]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 357.845 0.25 357.945 ;
			LAYER	M2 ;
			RECT	0 357.845 0.25 357.945 ;
			LAYER	M3 ;
			RECT	0 357.845 0.25 357.945 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[108]

	PIN DB[109]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 360.725 0.25 360.825 ;
			LAYER	M2 ;
			RECT	0 360.725 0.25 360.825 ;
			LAYER	M3 ;
			RECT	0 360.725 0.25 360.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[109]

	PIN DB[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 30.995 0.25 31.095 ;
			LAYER	M2 ;
			RECT	0 30.995 0.25 31.095 ;
			LAYER	M3 ;
			RECT	0 30.995 0.25 31.095 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[10]

	PIN DB[110]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 363.605 0.25 363.705 ;
			LAYER	M2 ;
			RECT	0 363.605 0.25 363.705 ;
			LAYER	M3 ;
			RECT	0 363.605 0.25 363.705 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[110]

	PIN DB[111]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 366.485 0.25 366.585 ;
			LAYER	M2 ;
			RECT	0 366.485 0.25 366.585 ;
			LAYER	M3 ;
			RECT	0 366.485 0.25 366.585 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[111]

	PIN DB[112]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 369.365 0.25 369.465 ;
			LAYER	M2 ;
			RECT	0 369.365 0.25 369.465 ;
			LAYER	M3 ;
			RECT	0 369.365 0.25 369.465 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[112]

	PIN DB[113]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 372.245 0.25 372.345 ;
			LAYER	M2 ;
			RECT	0 372.245 0.25 372.345 ;
			LAYER	M3 ;
			RECT	0 372.245 0.25 372.345 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[113]

	PIN DB[114]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 375.125 0.25 375.225 ;
			LAYER	M2 ;
			RECT	0 375.125 0.25 375.225 ;
			LAYER	M3 ;
			RECT	0 375.125 0.25 375.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[114]

	PIN DB[115]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 378.005 0.25 378.105 ;
			LAYER	M2 ;
			RECT	0 378.005 0.25 378.105 ;
			LAYER	M3 ;
			RECT	0 378.005 0.25 378.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[115]

	PIN DB[116]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 380.885 0.25 380.985 ;
			LAYER	M2 ;
			RECT	0 380.885 0.25 380.985 ;
			LAYER	M3 ;
			RECT	0 380.885 0.25 380.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[116]

	PIN DB[117]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 383.765 0.25 383.865 ;
			LAYER	M2 ;
			RECT	0 383.765 0.25 383.865 ;
			LAYER	M3 ;
			RECT	0 383.765 0.25 383.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[117]

	PIN DB[118]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 386.645 0.25 386.745 ;
			LAYER	M2 ;
			RECT	0 386.645 0.25 386.745 ;
			LAYER	M3 ;
			RECT	0 386.645 0.25 386.745 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[118]

	PIN DB[119]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 389.525 0.25 389.625 ;
			LAYER	M2 ;
			RECT	0 389.525 0.25 389.625 ;
			LAYER	M3 ;
			RECT	0 389.525 0.25 389.625 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[119]

	PIN DB[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 33.875 0.25 33.975 ;
			LAYER	M2 ;
			RECT	0 33.875 0.25 33.975 ;
			LAYER	M3 ;
			RECT	0 33.875 0.25 33.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[11]

	PIN DB[120]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 392.405 0.25 392.505 ;
			LAYER	M2 ;
			RECT	0 392.405 0.25 392.505 ;
			LAYER	M3 ;
			RECT	0 392.405 0.25 392.505 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[120]

	PIN DB[121]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 395.285 0.25 395.385 ;
			LAYER	M2 ;
			RECT	0 395.285 0.25 395.385 ;
			LAYER	M3 ;
			RECT	0 395.285 0.25 395.385 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[121]

	PIN DB[122]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 398.165 0.25 398.265 ;
			LAYER	M2 ;
			RECT	0 398.165 0.25 398.265 ;
			LAYER	M3 ;
			RECT	0 398.165 0.25 398.265 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[122]

	PIN DB[123]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 401.045 0.25 401.145 ;
			LAYER	M2 ;
			RECT	0 401.045 0.25 401.145 ;
			LAYER	M3 ;
			RECT	0 401.045 0.25 401.145 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[123]

	PIN DB[124]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 403.925 0.25 404.025 ;
			LAYER	M2 ;
			RECT	0 403.925 0.25 404.025 ;
			LAYER	M3 ;
			RECT	0 403.925 0.25 404.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[124]

	PIN DB[125]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 406.805 0.25 406.905 ;
			LAYER	M2 ;
			RECT	0 406.805 0.25 406.905 ;
			LAYER	M3 ;
			RECT	0 406.805 0.25 406.905 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[125]

	PIN DB[126]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 409.685 0.25 409.785 ;
			LAYER	M2 ;
			RECT	0 409.685 0.25 409.785 ;
			LAYER	M3 ;
			RECT	0 409.685 0.25 409.785 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[126]

	PIN DB[127]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 412.565 0.25 412.665 ;
			LAYER	M2 ;
			RECT	0 412.565 0.25 412.665 ;
			LAYER	M3 ;
			RECT	0 412.565 0.25 412.665 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[127]

	PIN DB[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 36.755 0.25 36.855 ;
			LAYER	M2 ;
			RECT	0 36.755 0.25 36.855 ;
			LAYER	M3 ;
			RECT	0 36.755 0.25 36.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[12]

	PIN DB[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 39.635 0.25 39.735 ;
			LAYER	M2 ;
			RECT	0 39.635 0.25 39.735 ;
			LAYER	M3 ;
			RECT	0 39.635 0.25 39.735 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[13]

	PIN DB[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 42.515 0.25 42.615 ;
			LAYER	M2 ;
			RECT	0 42.515 0.25 42.615 ;
			LAYER	M3 ;
			RECT	0 42.515 0.25 42.615 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[14]

	PIN DB[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 45.395 0.25 45.495 ;
			LAYER	M2 ;
			RECT	0 45.395 0.25 45.495 ;
			LAYER	M3 ;
			RECT	0 45.395 0.25 45.495 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[15]

	PIN DB[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 48.275 0.25 48.375 ;
			LAYER	M2 ;
			RECT	0 48.275 0.25 48.375 ;
			LAYER	M3 ;
			RECT	0 48.275 0.25 48.375 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[16]

	PIN DB[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 51.155 0.25 51.255 ;
			LAYER	M2 ;
			RECT	0 51.155 0.25 51.255 ;
			LAYER	M3 ;
			RECT	0 51.155 0.25 51.255 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[17]

	PIN DB[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 54.035 0.25 54.135 ;
			LAYER	M2 ;
			RECT	0 54.035 0.25 54.135 ;
			LAYER	M3 ;
			RECT	0 54.035 0.25 54.135 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[18]

	PIN DB[19]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 56.915 0.25 57.015 ;
			LAYER	M2 ;
			RECT	0 56.915 0.25 57.015 ;
			LAYER	M3 ;
			RECT	0 56.915 0.25 57.015 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[19]

	PIN DB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 5.075 0.25 5.175 ;
			LAYER	M2 ;
			RECT	0 5.075 0.25 5.175 ;
			LAYER	M3 ;
			RECT	0 5.075 0.25 5.175 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[1]

	PIN DB[20]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 59.795 0.25 59.895 ;
			LAYER	M2 ;
			RECT	0 59.795 0.25 59.895 ;
			LAYER	M3 ;
			RECT	0 59.795 0.25 59.895 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[20]

	PIN DB[21]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 62.675 0.25 62.775 ;
			LAYER	M2 ;
			RECT	0 62.675 0.25 62.775 ;
			LAYER	M3 ;
			RECT	0 62.675 0.25 62.775 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[21]

	PIN DB[22]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 65.555 0.25 65.655 ;
			LAYER	M2 ;
			RECT	0 65.555 0.25 65.655 ;
			LAYER	M3 ;
			RECT	0 65.555 0.25 65.655 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[22]

	PIN DB[23]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 68.435 0.25 68.535 ;
			LAYER	M2 ;
			RECT	0 68.435 0.25 68.535 ;
			LAYER	M3 ;
			RECT	0 68.435 0.25 68.535 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[23]

	PIN DB[24]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 71.315 0.25 71.415 ;
			LAYER	M2 ;
			RECT	0 71.315 0.25 71.415 ;
			LAYER	M3 ;
			RECT	0 71.315 0.25 71.415 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[24]

	PIN DB[25]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 74.195 0.25 74.295 ;
			LAYER	M2 ;
			RECT	0 74.195 0.25 74.295 ;
			LAYER	M3 ;
			RECT	0 74.195 0.25 74.295 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[25]

	PIN DB[26]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 77.075 0.25 77.175 ;
			LAYER	M2 ;
			RECT	0 77.075 0.25 77.175 ;
			LAYER	M3 ;
			RECT	0 77.075 0.25 77.175 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[26]

	PIN DB[27]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 79.955 0.25 80.055 ;
			LAYER	M2 ;
			RECT	0 79.955 0.25 80.055 ;
			LAYER	M3 ;
			RECT	0 79.955 0.25 80.055 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[27]

	PIN DB[28]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 82.835 0.25 82.935 ;
			LAYER	M2 ;
			RECT	0 82.835 0.25 82.935 ;
			LAYER	M3 ;
			RECT	0 82.835 0.25 82.935 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[28]

	PIN DB[29]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 85.715 0.25 85.815 ;
			LAYER	M2 ;
			RECT	0 85.715 0.25 85.815 ;
			LAYER	M3 ;
			RECT	0 85.715 0.25 85.815 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[29]

	PIN DB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 7.955 0.25 8.055 ;
			LAYER	M2 ;
			RECT	0 7.955 0.25 8.055 ;
			LAYER	M3 ;
			RECT	0 7.955 0.25 8.055 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[2]

	PIN DB[30]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 88.595 0.25 88.695 ;
			LAYER	M2 ;
			RECT	0 88.595 0.25 88.695 ;
			LAYER	M3 ;
			RECT	0 88.595 0.25 88.695 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[30]

	PIN DB[31]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 91.475 0.25 91.575 ;
			LAYER	M2 ;
			RECT	0 91.475 0.25 91.575 ;
			LAYER	M3 ;
			RECT	0 91.475 0.25 91.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[31]

	PIN DB[32]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 94.355 0.25 94.455 ;
			LAYER	M2 ;
			RECT	0 94.355 0.25 94.455 ;
			LAYER	M3 ;
			RECT	0 94.355 0.25 94.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[32]

	PIN DB[33]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 97.235 0.25 97.335 ;
			LAYER	M2 ;
			RECT	0 97.235 0.25 97.335 ;
			LAYER	M3 ;
			RECT	0 97.235 0.25 97.335 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[33]

	PIN DB[34]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 100.115 0.25 100.215 ;
			LAYER	M2 ;
			RECT	0 100.115 0.25 100.215 ;
			LAYER	M3 ;
			RECT	0 100.115 0.25 100.215 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[34]

	PIN DB[35]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 102.995 0.25 103.095 ;
			LAYER	M2 ;
			RECT	0 102.995 0.25 103.095 ;
			LAYER	M3 ;
			RECT	0 102.995 0.25 103.095 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[35]

	PIN DB[36]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 105.875 0.25 105.975 ;
			LAYER	M2 ;
			RECT	0 105.875 0.25 105.975 ;
			LAYER	M3 ;
			RECT	0 105.875 0.25 105.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[36]

	PIN DB[37]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 108.755 0.25 108.855 ;
			LAYER	M2 ;
			RECT	0 108.755 0.25 108.855 ;
			LAYER	M3 ;
			RECT	0 108.755 0.25 108.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[37]

	PIN DB[38]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 111.635 0.25 111.735 ;
			LAYER	M2 ;
			RECT	0 111.635 0.25 111.735 ;
			LAYER	M3 ;
			RECT	0 111.635 0.25 111.735 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[38]

	PIN DB[39]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 114.515 0.25 114.615 ;
			LAYER	M2 ;
			RECT	0 114.515 0.25 114.615 ;
			LAYER	M3 ;
			RECT	0 114.515 0.25 114.615 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[39]

	PIN DB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 10.835 0.25 10.935 ;
			LAYER	M2 ;
			RECT	0 10.835 0.25 10.935 ;
			LAYER	M3 ;
			RECT	0 10.835 0.25 10.935 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[3]

	PIN DB[40]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 117.395 0.25 117.495 ;
			LAYER	M2 ;
			RECT	0 117.395 0.25 117.495 ;
			LAYER	M3 ;
			RECT	0 117.395 0.25 117.495 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[40]

	PIN DB[41]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 120.275 0.25 120.375 ;
			LAYER	M2 ;
			RECT	0 120.275 0.25 120.375 ;
			LAYER	M3 ;
			RECT	0 120.275 0.25 120.375 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[41]

	PIN DB[42]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 123.155 0.25 123.255 ;
			LAYER	M2 ;
			RECT	0 123.155 0.25 123.255 ;
			LAYER	M3 ;
			RECT	0 123.155 0.25 123.255 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[42]

	PIN DB[43]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 126.035 0.25 126.135 ;
			LAYER	M2 ;
			RECT	0 126.035 0.25 126.135 ;
			LAYER	M3 ;
			RECT	0 126.035 0.25 126.135 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[43]

	PIN DB[44]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 128.915 0.25 129.015 ;
			LAYER	M2 ;
			RECT	0 128.915 0.25 129.015 ;
			LAYER	M3 ;
			RECT	0 128.915 0.25 129.015 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[44]

	PIN DB[45]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 131.795 0.25 131.895 ;
			LAYER	M2 ;
			RECT	0 131.795 0.25 131.895 ;
			LAYER	M3 ;
			RECT	0 131.795 0.25 131.895 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[45]

	PIN DB[46]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 134.675 0.25 134.775 ;
			LAYER	M2 ;
			RECT	0 134.675 0.25 134.775 ;
			LAYER	M3 ;
			RECT	0 134.675 0.25 134.775 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[46]

	PIN DB[47]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 137.555 0.25 137.655 ;
			LAYER	M2 ;
			RECT	0 137.555 0.25 137.655 ;
			LAYER	M3 ;
			RECT	0 137.555 0.25 137.655 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[47]

	PIN DB[48]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 140.435 0.25 140.535 ;
			LAYER	M2 ;
			RECT	0 140.435 0.25 140.535 ;
			LAYER	M3 ;
			RECT	0 140.435 0.25 140.535 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[48]

	PIN DB[49]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 143.315 0.25 143.415 ;
			LAYER	M2 ;
			RECT	0 143.315 0.25 143.415 ;
			LAYER	M3 ;
			RECT	0 143.315 0.25 143.415 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[49]

	PIN DB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 13.715 0.25 13.815 ;
			LAYER	M2 ;
			RECT	0 13.715 0.25 13.815 ;
			LAYER	M3 ;
			RECT	0 13.715 0.25 13.815 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[4]

	PIN DB[50]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 146.195 0.25 146.295 ;
			LAYER	M2 ;
			RECT	0 146.195 0.25 146.295 ;
			LAYER	M3 ;
			RECT	0 146.195 0.25 146.295 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[50]

	PIN DB[51]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 149.075 0.25 149.175 ;
			LAYER	M2 ;
			RECT	0 149.075 0.25 149.175 ;
			LAYER	M3 ;
			RECT	0 149.075 0.25 149.175 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[51]

	PIN DB[52]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 151.955 0.25 152.055 ;
			LAYER	M2 ;
			RECT	0 151.955 0.25 152.055 ;
			LAYER	M3 ;
			RECT	0 151.955 0.25 152.055 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[52]

	PIN DB[53]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 154.835 0.25 154.935 ;
			LAYER	M2 ;
			RECT	0 154.835 0.25 154.935 ;
			LAYER	M3 ;
			RECT	0 154.835 0.25 154.935 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[53]

	PIN DB[54]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 157.715 0.25 157.815 ;
			LAYER	M2 ;
			RECT	0 157.715 0.25 157.815 ;
			LAYER	M3 ;
			RECT	0 157.715 0.25 157.815 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[54]

	PIN DB[55]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 160.595 0.25 160.695 ;
			LAYER	M2 ;
			RECT	0 160.595 0.25 160.695 ;
			LAYER	M3 ;
			RECT	0 160.595 0.25 160.695 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[55]

	PIN DB[56]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 163.475 0.25 163.575 ;
			LAYER	M2 ;
			RECT	0 163.475 0.25 163.575 ;
			LAYER	M3 ;
			RECT	0 163.475 0.25 163.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[56]

	PIN DB[57]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 166.355 0.25 166.455 ;
			LAYER	M2 ;
			RECT	0 166.355 0.25 166.455 ;
			LAYER	M3 ;
			RECT	0 166.355 0.25 166.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[57]

	PIN DB[58]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 169.235 0.25 169.335 ;
			LAYER	M2 ;
			RECT	0 169.235 0.25 169.335 ;
			LAYER	M3 ;
			RECT	0 169.235 0.25 169.335 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[58]

	PIN DB[59]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 172.115 0.25 172.215 ;
			LAYER	M2 ;
			RECT	0 172.115 0.25 172.215 ;
			LAYER	M3 ;
			RECT	0 172.115 0.25 172.215 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[59]

	PIN DB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 16.595 0.25 16.695 ;
			LAYER	M2 ;
			RECT	0 16.595 0.25 16.695 ;
			LAYER	M3 ;
			RECT	0 16.595 0.25 16.695 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[5]

	PIN DB[60]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 174.995 0.25 175.095 ;
			LAYER	M2 ;
			RECT	0 174.995 0.25 175.095 ;
			LAYER	M3 ;
			RECT	0 174.995 0.25 175.095 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[60]

	PIN DB[61]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 177.875 0.25 177.975 ;
			LAYER	M2 ;
			RECT	0 177.875 0.25 177.975 ;
			LAYER	M3 ;
			RECT	0 177.875 0.25 177.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[61]

	PIN DB[62]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 180.755 0.25 180.855 ;
			LAYER	M2 ;
			RECT	0 180.755 0.25 180.855 ;
			LAYER	M3 ;
			RECT	0 180.755 0.25 180.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[62]

	PIN DB[63]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 183.635 0.25 183.735 ;
			LAYER	M2 ;
			RECT	0 183.635 0.25 183.735 ;
			LAYER	M3 ;
			RECT	0 183.635 0.25 183.735 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[63]

	PIN DB[64]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 231.125 0.25 231.225 ;
			LAYER	M2 ;
			RECT	0 231.125 0.25 231.225 ;
			LAYER	M3 ;
			RECT	0 231.125 0.25 231.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[64]

	PIN DB[65]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 234.005 0.25 234.105 ;
			LAYER	M2 ;
			RECT	0 234.005 0.25 234.105 ;
			LAYER	M3 ;
			RECT	0 234.005 0.25 234.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[65]

	PIN DB[66]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 236.885 0.25 236.985 ;
			LAYER	M2 ;
			RECT	0 236.885 0.25 236.985 ;
			LAYER	M3 ;
			RECT	0 236.885 0.25 236.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[66]

	PIN DB[67]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 239.765 0.25 239.865 ;
			LAYER	M2 ;
			RECT	0 239.765 0.25 239.865 ;
			LAYER	M3 ;
			RECT	0 239.765 0.25 239.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[67]

	PIN DB[68]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 242.645 0.25 242.745 ;
			LAYER	M2 ;
			RECT	0 242.645 0.25 242.745 ;
			LAYER	M3 ;
			RECT	0 242.645 0.25 242.745 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[68]

	PIN DB[69]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 245.525 0.25 245.625 ;
			LAYER	M2 ;
			RECT	0 245.525 0.25 245.625 ;
			LAYER	M3 ;
			RECT	0 245.525 0.25 245.625 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[69]

	PIN DB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 19.475 0.25 19.575 ;
			LAYER	M2 ;
			RECT	0 19.475 0.25 19.575 ;
			LAYER	M3 ;
			RECT	0 19.475 0.25 19.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[6]

	PIN DB[70]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 248.405 0.25 248.505 ;
			LAYER	M2 ;
			RECT	0 248.405 0.25 248.505 ;
			LAYER	M3 ;
			RECT	0 248.405 0.25 248.505 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[70]

	PIN DB[71]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 251.285 0.25 251.385 ;
			LAYER	M2 ;
			RECT	0 251.285 0.25 251.385 ;
			LAYER	M3 ;
			RECT	0 251.285 0.25 251.385 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[71]

	PIN DB[72]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 254.165 0.25 254.265 ;
			LAYER	M2 ;
			RECT	0 254.165 0.25 254.265 ;
			LAYER	M3 ;
			RECT	0 254.165 0.25 254.265 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[72]

	PIN DB[73]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 257.045 0.25 257.145 ;
			LAYER	M2 ;
			RECT	0 257.045 0.25 257.145 ;
			LAYER	M3 ;
			RECT	0 257.045 0.25 257.145 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[73]

	PIN DB[74]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 259.925 0.25 260.025 ;
			LAYER	M2 ;
			RECT	0 259.925 0.25 260.025 ;
			LAYER	M3 ;
			RECT	0 259.925 0.25 260.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[74]

	PIN DB[75]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 262.805 0.25 262.905 ;
			LAYER	M2 ;
			RECT	0 262.805 0.25 262.905 ;
			LAYER	M3 ;
			RECT	0 262.805 0.25 262.905 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[75]

	PIN DB[76]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 265.685 0.25 265.785 ;
			LAYER	M2 ;
			RECT	0 265.685 0.25 265.785 ;
			LAYER	M3 ;
			RECT	0 265.685 0.25 265.785 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[76]

	PIN DB[77]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 268.565 0.25 268.665 ;
			LAYER	M2 ;
			RECT	0 268.565 0.25 268.665 ;
			LAYER	M3 ;
			RECT	0 268.565 0.25 268.665 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[77]

	PIN DB[78]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 271.445 0.25 271.545 ;
			LAYER	M2 ;
			RECT	0 271.445 0.25 271.545 ;
			LAYER	M3 ;
			RECT	0 271.445 0.25 271.545 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[78]

	PIN DB[79]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 274.325 0.25 274.425 ;
			LAYER	M2 ;
			RECT	0 274.325 0.25 274.425 ;
			LAYER	M3 ;
			RECT	0 274.325 0.25 274.425 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[79]

	PIN DB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 22.355 0.25 22.455 ;
			LAYER	M2 ;
			RECT	0 22.355 0.25 22.455 ;
			LAYER	M3 ;
			RECT	0 22.355 0.25 22.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[7]

	PIN DB[80]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 277.205 0.25 277.305 ;
			LAYER	M2 ;
			RECT	0 277.205 0.25 277.305 ;
			LAYER	M3 ;
			RECT	0 277.205 0.25 277.305 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[80]

	PIN DB[81]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 280.085 0.25 280.185 ;
			LAYER	M2 ;
			RECT	0 280.085 0.25 280.185 ;
			LAYER	M3 ;
			RECT	0 280.085 0.25 280.185 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[81]

	PIN DB[82]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 282.965 0.25 283.065 ;
			LAYER	M2 ;
			RECT	0 282.965 0.25 283.065 ;
			LAYER	M3 ;
			RECT	0 282.965 0.25 283.065 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[82]

	PIN DB[83]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 285.845 0.25 285.945 ;
			LAYER	M2 ;
			RECT	0 285.845 0.25 285.945 ;
			LAYER	M3 ;
			RECT	0 285.845 0.25 285.945 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[83]

	PIN DB[84]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 288.725 0.25 288.825 ;
			LAYER	M2 ;
			RECT	0 288.725 0.25 288.825 ;
			LAYER	M3 ;
			RECT	0 288.725 0.25 288.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[84]

	PIN DB[85]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 291.605 0.25 291.705 ;
			LAYER	M2 ;
			RECT	0 291.605 0.25 291.705 ;
			LAYER	M3 ;
			RECT	0 291.605 0.25 291.705 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[85]

	PIN DB[86]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 294.485 0.25 294.585 ;
			LAYER	M2 ;
			RECT	0 294.485 0.25 294.585 ;
			LAYER	M3 ;
			RECT	0 294.485 0.25 294.585 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[86]

	PIN DB[87]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 297.365 0.25 297.465 ;
			LAYER	M2 ;
			RECT	0 297.365 0.25 297.465 ;
			LAYER	M3 ;
			RECT	0 297.365 0.25 297.465 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[87]

	PIN DB[88]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 300.245 0.25 300.345 ;
			LAYER	M2 ;
			RECT	0 300.245 0.25 300.345 ;
			LAYER	M3 ;
			RECT	0 300.245 0.25 300.345 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[88]

	PIN DB[89]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 303.125 0.25 303.225 ;
			LAYER	M2 ;
			RECT	0 303.125 0.25 303.225 ;
			LAYER	M3 ;
			RECT	0 303.125 0.25 303.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[89]

	PIN DB[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 25.235 0.25 25.335 ;
			LAYER	M2 ;
			RECT	0 25.235 0.25 25.335 ;
			LAYER	M3 ;
			RECT	0 25.235 0.25 25.335 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[8]

	PIN DB[90]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 306.005 0.25 306.105 ;
			LAYER	M2 ;
			RECT	0 306.005 0.25 306.105 ;
			LAYER	M3 ;
			RECT	0 306.005 0.25 306.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[90]

	PIN DB[91]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 308.885 0.25 308.985 ;
			LAYER	M2 ;
			RECT	0 308.885 0.25 308.985 ;
			LAYER	M3 ;
			RECT	0 308.885 0.25 308.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[91]

	PIN DB[92]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 311.765 0.25 311.865 ;
			LAYER	M2 ;
			RECT	0 311.765 0.25 311.865 ;
			LAYER	M3 ;
			RECT	0 311.765 0.25 311.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[92]

	PIN DB[93]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 314.645 0.25 314.745 ;
			LAYER	M2 ;
			RECT	0 314.645 0.25 314.745 ;
			LAYER	M3 ;
			RECT	0 314.645 0.25 314.745 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[93]

	PIN DB[94]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 317.525 0.25 317.625 ;
			LAYER	M2 ;
			RECT	0 317.525 0.25 317.625 ;
			LAYER	M3 ;
			RECT	0 317.525 0.25 317.625 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[94]

	PIN DB[95]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 320.405 0.25 320.505 ;
			LAYER	M2 ;
			RECT	0 320.405 0.25 320.505 ;
			LAYER	M3 ;
			RECT	0 320.405 0.25 320.505 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[95]

	PIN DB[96]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 323.285 0.25 323.385 ;
			LAYER	M2 ;
			RECT	0 323.285 0.25 323.385 ;
			LAYER	M3 ;
			RECT	0 323.285 0.25 323.385 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[96]

	PIN DB[97]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 326.165 0.25 326.265 ;
			LAYER	M2 ;
			RECT	0 326.165 0.25 326.265 ;
			LAYER	M3 ;
			RECT	0 326.165 0.25 326.265 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[97]

	PIN DB[98]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 329.045 0.25 329.145 ;
			LAYER	M2 ;
			RECT	0 329.045 0.25 329.145 ;
			LAYER	M3 ;
			RECT	0 329.045 0.25 329.145 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[98]

	PIN DB[99]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 331.925 0.25 332.025 ;
			LAYER	M2 ;
			RECT	0 331.925 0.25 332.025 ;
			LAYER	M3 ;
			RECT	0 331.925 0.25 332.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[99]

	PIN DB[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 28.115 0.25 28.215 ;
			LAYER	M2 ;
			RECT	0 28.115 0.25 28.215 ;
			LAYER	M3 ;
			RECT	0 28.115 0.25 28.215 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[9]

	PIN DFTRAMBYP
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 225.7 0.25 225.8 ;
			LAYER	M2 ;
			RECT	0 225.7 0.25 225.8 ;
			LAYER	M3 ;
			RECT	0 225.7 0.25 225.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DFTRAMBYP

	PIN EMAA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 199.77 0.25 199.87 ;
			LAYER	M2 ;
			RECT	0 199.77 0.25 199.87 ;
			LAYER	M3 ;
			RECT	0 199.77 0.25 199.87 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAA[0]

	PIN EMAA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 199.57 0.25 199.67 ;
			LAYER	M2 ;
			RECT	0 199.57 0.25 199.67 ;
			LAYER	M3 ;
			RECT	0 199.57 0.25 199.67 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAA[1]

	PIN EMAA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 201.505 0.25 201.605 ;
			LAYER	M2 ;
			RECT	0 201.505 0.25 201.605 ;
			LAYER	M3 ;
			RECT	0 201.505 0.25 201.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAA[2]

	PIN EMAB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 214.305 0.25 214.405 ;
			LAYER	M2 ;
			RECT	0 214.305 0.25 214.405 ;
			LAYER	M3 ;
			RECT	0 214.305 0.25 214.405 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAB[0]

	PIN EMAB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 215.305 0.25 215.405 ;
			LAYER	M2 ;
			RECT	0 215.305 0.25 215.405 ;
			LAYER	M3 ;
			RECT	0 215.305 0.25 215.405 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAB[1]

	PIN EMAB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 212.825 0.25 212.925 ;
			LAYER	M2 ;
			RECT	0 212.825 0.25 212.925 ;
			LAYER	M3 ;
			RECT	0 212.825 0.25 212.925 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAB[2]

	PIN EMASA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 187.45 0.25 187.55 ;
			LAYER	M2 ;
			RECT	0 187.45 0.25 187.55 ;
			LAYER	M3 ;
			RECT	0 187.45 0.25 187.55 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMASA

	PIN QA[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 2.455 0.25 2.555 ;
			LAYER	M2 ;
			RECT	0 2.455 0.25 2.555 ;
			LAYER	M3 ;
			RECT	0 2.455 0.25 2.555 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[0]

	PIN QA[100]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 334.545 0.25 334.645 ;
			LAYER	M2 ;
			RECT	0 334.545 0.25 334.645 ;
			LAYER	M3 ;
			RECT	0 334.545 0.25 334.645 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[100]

	PIN QA[101]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 337.425 0.25 337.525 ;
			LAYER	M2 ;
			RECT	0 337.425 0.25 337.525 ;
			LAYER	M3 ;
			RECT	0 337.425 0.25 337.525 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[101]

	PIN QA[102]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 340.305 0.25 340.405 ;
			LAYER	M2 ;
			RECT	0 340.305 0.25 340.405 ;
			LAYER	M3 ;
			RECT	0 340.305 0.25 340.405 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[102]

	PIN QA[103]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 343.185 0.25 343.285 ;
			LAYER	M2 ;
			RECT	0 343.185 0.25 343.285 ;
			LAYER	M3 ;
			RECT	0 343.185 0.25 343.285 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[103]

	PIN QA[104]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 346.065 0.25 346.165 ;
			LAYER	M2 ;
			RECT	0 346.065 0.25 346.165 ;
			LAYER	M3 ;
			RECT	0 346.065 0.25 346.165 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[104]

	PIN QA[105]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 348.945 0.25 349.045 ;
			LAYER	M2 ;
			RECT	0 348.945 0.25 349.045 ;
			LAYER	M3 ;
			RECT	0 348.945 0.25 349.045 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[105]

	PIN QA[106]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 351.825 0.25 351.925 ;
			LAYER	M2 ;
			RECT	0 351.825 0.25 351.925 ;
			LAYER	M3 ;
			RECT	0 351.825 0.25 351.925 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[106]

	PIN QA[107]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 354.705 0.25 354.805 ;
			LAYER	M2 ;
			RECT	0 354.705 0.25 354.805 ;
			LAYER	M3 ;
			RECT	0 354.705 0.25 354.805 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[107]

	PIN QA[108]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 357.585 0.25 357.685 ;
			LAYER	M2 ;
			RECT	0 357.585 0.25 357.685 ;
			LAYER	M3 ;
			RECT	0 357.585 0.25 357.685 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[108]

	PIN QA[109]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 360.465 0.25 360.565 ;
			LAYER	M2 ;
			RECT	0 360.465 0.25 360.565 ;
			LAYER	M3 ;
			RECT	0 360.465 0.25 360.565 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[109]

	PIN QA[10]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 31.255 0.25 31.355 ;
			LAYER	M2 ;
			RECT	0 31.255 0.25 31.355 ;
			LAYER	M3 ;
			RECT	0 31.255 0.25 31.355 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[10]

	PIN QA[110]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 363.345 0.25 363.445 ;
			LAYER	M2 ;
			RECT	0 363.345 0.25 363.445 ;
			LAYER	M3 ;
			RECT	0 363.345 0.25 363.445 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[110]

	PIN QA[111]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 366.225 0.25 366.325 ;
			LAYER	M2 ;
			RECT	0 366.225 0.25 366.325 ;
			LAYER	M3 ;
			RECT	0 366.225 0.25 366.325 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[111]

	PIN QA[112]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 369.105 0.25 369.205 ;
			LAYER	M2 ;
			RECT	0 369.105 0.25 369.205 ;
			LAYER	M3 ;
			RECT	0 369.105 0.25 369.205 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[112]

	PIN QA[113]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 371.985 0.25 372.085 ;
			LAYER	M2 ;
			RECT	0 371.985 0.25 372.085 ;
			LAYER	M3 ;
			RECT	0 371.985 0.25 372.085 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[113]

	PIN QA[114]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 374.865 0.25 374.965 ;
			LAYER	M2 ;
			RECT	0 374.865 0.25 374.965 ;
			LAYER	M3 ;
			RECT	0 374.865 0.25 374.965 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[114]

	PIN QA[115]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 377.745 0.25 377.845 ;
			LAYER	M2 ;
			RECT	0 377.745 0.25 377.845 ;
			LAYER	M3 ;
			RECT	0 377.745 0.25 377.845 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[115]

	PIN QA[116]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 380.625 0.25 380.725 ;
			LAYER	M2 ;
			RECT	0 380.625 0.25 380.725 ;
			LAYER	M3 ;
			RECT	0 380.625 0.25 380.725 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[116]

	PIN QA[117]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 383.505 0.25 383.605 ;
			LAYER	M2 ;
			RECT	0 383.505 0.25 383.605 ;
			LAYER	M3 ;
			RECT	0 383.505 0.25 383.605 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[117]

	PIN QA[118]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 386.385 0.25 386.485 ;
			LAYER	M2 ;
			RECT	0 386.385 0.25 386.485 ;
			LAYER	M3 ;
			RECT	0 386.385 0.25 386.485 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[118]

	PIN QA[119]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 389.265 0.25 389.365 ;
			LAYER	M2 ;
			RECT	0 389.265 0.25 389.365 ;
			LAYER	M3 ;
			RECT	0 389.265 0.25 389.365 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[119]

	PIN QA[11]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 34.135 0.25 34.235 ;
			LAYER	M2 ;
			RECT	0 34.135 0.25 34.235 ;
			LAYER	M3 ;
			RECT	0 34.135 0.25 34.235 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[11]

	PIN QA[120]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 392.145 0.25 392.245 ;
			LAYER	M2 ;
			RECT	0 392.145 0.25 392.245 ;
			LAYER	M3 ;
			RECT	0 392.145 0.25 392.245 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[120]

	PIN QA[121]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 395.025 0.25 395.125 ;
			LAYER	M2 ;
			RECT	0 395.025 0.25 395.125 ;
			LAYER	M3 ;
			RECT	0 395.025 0.25 395.125 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[121]

	PIN QA[122]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 397.905 0.25 398.005 ;
			LAYER	M2 ;
			RECT	0 397.905 0.25 398.005 ;
			LAYER	M3 ;
			RECT	0 397.905 0.25 398.005 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[122]

	PIN QA[123]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 400.785 0.25 400.885 ;
			LAYER	M2 ;
			RECT	0 400.785 0.25 400.885 ;
			LAYER	M3 ;
			RECT	0 400.785 0.25 400.885 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[123]

	PIN QA[124]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 403.665 0.25 403.765 ;
			LAYER	M2 ;
			RECT	0 403.665 0.25 403.765 ;
			LAYER	M3 ;
			RECT	0 403.665 0.25 403.765 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[124]

	PIN QA[125]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 406.545 0.25 406.645 ;
			LAYER	M2 ;
			RECT	0 406.545 0.25 406.645 ;
			LAYER	M3 ;
			RECT	0 406.545 0.25 406.645 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[125]

	PIN QA[126]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 409.425 0.25 409.525 ;
			LAYER	M2 ;
			RECT	0 409.425 0.25 409.525 ;
			LAYER	M3 ;
			RECT	0 409.425 0.25 409.525 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[126]

	PIN QA[127]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 412.305 0.25 412.405 ;
			LAYER	M2 ;
			RECT	0 412.305 0.25 412.405 ;
			LAYER	M3 ;
			RECT	0 412.305 0.25 412.405 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[127]

	PIN QA[12]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 37.015 0.25 37.115 ;
			LAYER	M2 ;
			RECT	0 37.015 0.25 37.115 ;
			LAYER	M3 ;
			RECT	0 37.015 0.25 37.115 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[12]

	PIN QA[13]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 39.895 0.25 39.995 ;
			LAYER	M2 ;
			RECT	0 39.895 0.25 39.995 ;
			LAYER	M3 ;
			RECT	0 39.895 0.25 39.995 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[13]

	PIN QA[14]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 42.775 0.25 42.875 ;
			LAYER	M2 ;
			RECT	0 42.775 0.25 42.875 ;
			LAYER	M3 ;
			RECT	0 42.775 0.25 42.875 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[14]

	PIN QA[15]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 45.655 0.25 45.755 ;
			LAYER	M2 ;
			RECT	0 45.655 0.25 45.755 ;
			LAYER	M3 ;
			RECT	0 45.655 0.25 45.755 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[15]

	PIN QA[16]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 48.535 0.25 48.635 ;
			LAYER	M2 ;
			RECT	0 48.535 0.25 48.635 ;
			LAYER	M3 ;
			RECT	0 48.535 0.25 48.635 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[16]

	PIN QA[17]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 51.415 0.25 51.515 ;
			LAYER	M2 ;
			RECT	0 51.415 0.25 51.515 ;
			LAYER	M3 ;
			RECT	0 51.415 0.25 51.515 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[17]

	PIN QA[18]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 54.295 0.25 54.395 ;
			LAYER	M2 ;
			RECT	0 54.295 0.25 54.395 ;
			LAYER	M3 ;
			RECT	0 54.295 0.25 54.395 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[18]

	PIN QA[19]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 57.175 0.25 57.275 ;
			LAYER	M2 ;
			RECT	0 57.175 0.25 57.275 ;
			LAYER	M3 ;
			RECT	0 57.175 0.25 57.275 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[19]

	PIN QA[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 5.335 0.25 5.435 ;
			LAYER	M2 ;
			RECT	0 5.335 0.25 5.435 ;
			LAYER	M3 ;
			RECT	0 5.335 0.25 5.435 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[1]

	PIN QA[20]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 60.055 0.25 60.155 ;
			LAYER	M2 ;
			RECT	0 60.055 0.25 60.155 ;
			LAYER	M3 ;
			RECT	0 60.055 0.25 60.155 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[20]

	PIN QA[21]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 62.935 0.25 63.035 ;
			LAYER	M2 ;
			RECT	0 62.935 0.25 63.035 ;
			LAYER	M3 ;
			RECT	0 62.935 0.25 63.035 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[21]

	PIN QA[22]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 65.815 0.25 65.915 ;
			LAYER	M2 ;
			RECT	0 65.815 0.25 65.915 ;
			LAYER	M3 ;
			RECT	0 65.815 0.25 65.915 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[22]

	PIN QA[23]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 68.695 0.25 68.795 ;
			LAYER	M2 ;
			RECT	0 68.695 0.25 68.795 ;
			LAYER	M3 ;
			RECT	0 68.695 0.25 68.795 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[23]

	PIN QA[24]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 71.575 0.25 71.675 ;
			LAYER	M2 ;
			RECT	0 71.575 0.25 71.675 ;
			LAYER	M3 ;
			RECT	0 71.575 0.25 71.675 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[24]

	PIN QA[25]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 74.455 0.25 74.555 ;
			LAYER	M2 ;
			RECT	0 74.455 0.25 74.555 ;
			LAYER	M3 ;
			RECT	0 74.455 0.25 74.555 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[25]

	PIN QA[26]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 77.335 0.25 77.435 ;
			LAYER	M2 ;
			RECT	0 77.335 0.25 77.435 ;
			LAYER	M3 ;
			RECT	0 77.335 0.25 77.435 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[26]

	PIN QA[27]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 80.215 0.25 80.315 ;
			LAYER	M2 ;
			RECT	0 80.215 0.25 80.315 ;
			LAYER	M3 ;
			RECT	0 80.215 0.25 80.315 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[27]

	PIN QA[28]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 83.095 0.25 83.195 ;
			LAYER	M2 ;
			RECT	0 83.095 0.25 83.195 ;
			LAYER	M3 ;
			RECT	0 83.095 0.25 83.195 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[28]

	PIN QA[29]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 85.975 0.25 86.075 ;
			LAYER	M2 ;
			RECT	0 85.975 0.25 86.075 ;
			LAYER	M3 ;
			RECT	0 85.975 0.25 86.075 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[29]

	PIN QA[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 8.215 0.25 8.315 ;
			LAYER	M2 ;
			RECT	0 8.215 0.25 8.315 ;
			LAYER	M3 ;
			RECT	0 8.215 0.25 8.315 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[2]

	PIN QA[30]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 88.855 0.25 88.955 ;
			LAYER	M2 ;
			RECT	0 88.855 0.25 88.955 ;
			LAYER	M3 ;
			RECT	0 88.855 0.25 88.955 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[30]

	PIN QA[31]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 91.735 0.25 91.835 ;
			LAYER	M2 ;
			RECT	0 91.735 0.25 91.835 ;
			LAYER	M3 ;
			RECT	0 91.735 0.25 91.835 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[31]

	PIN QA[32]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 94.615 0.25 94.715 ;
			LAYER	M2 ;
			RECT	0 94.615 0.25 94.715 ;
			LAYER	M3 ;
			RECT	0 94.615 0.25 94.715 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[32]

	PIN QA[33]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 97.495 0.25 97.595 ;
			LAYER	M2 ;
			RECT	0 97.495 0.25 97.595 ;
			LAYER	M3 ;
			RECT	0 97.495 0.25 97.595 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[33]

	PIN QA[34]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 100.375 0.25 100.475 ;
			LAYER	M2 ;
			RECT	0 100.375 0.25 100.475 ;
			LAYER	M3 ;
			RECT	0 100.375 0.25 100.475 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[34]

	PIN QA[35]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 103.255 0.25 103.355 ;
			LAYER	M2 ;
			RECT	0 103.255 0.25 103.355 ;
			LAYER	M3 ;
			RECT	0 103.255 0.25 103.355 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[35]

	PIN QA[36]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 106.135 0.25 106.235 ;
			LAYER	M2 ;
			RECT	0 106.135 0.25 106.235 ;
			LAYER	M3 ;
			RECT	0 106.135 0.25 106.235 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[36]

	PIN QA[37]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 109.015 0.25 109.115 ;
			LAYER	M2 ;
			RECT	0 109.015 0.25 109.115 ;
			LAYER	M3 ;
			RECT	0 109.015 0.25 109.115 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[37]

	PIN QA[38]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 111.895 0.25 111.995 ;
			LAYER	M2 ;
			RECT	0 111.895 0.25 111.995 ;
			LAYER	M3 ;
			RECT	0 111.895 0.25 111.995 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[38]

	PIN QA[39]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 114.775 0.25 114.875 ;
			LAYER	M2 ;
			RECT	0 114.775 0.25 114.875 ;
			LAYER	M3 ;
			RECT	0 114.775 0.25 114.875 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[39]

	PIN QA[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 11.095 0.25 11.195 ;
			LAYER	M2 ;
			RECT	0 11.095 0.25 11.195 ;
			LAYER	M3 ;
			RECT	0 11.095 0.25 11.195 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[3]

	PIN QA[40]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 117.655 0.25 117.755 ;
			LAYER	M2 ;
			RECT	0 117.655 0.25 117.755 ;
			LAYER	M3 ;
			RECT	0 117.655 0.25 117.755 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[40]

	PIN QA[41]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 120.535 0.25 120.635 ;
			LAYER	M2 ;
			RECT	0 120.535 0.25 120.635 ;
			LAYER	M3 ;
			RECT	0 120.535 0.25 120.635 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[41]

	PIN QA[42]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 123.415 0.25 123.515 ;
			LAYER	M2 ;
			RECT	0 123.415 0.25 123.515 ;
			LAYER	M3 ;
			RECT	0 123.415 0.25 123.515 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[42]

	PIN QA[43]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 126.295 0.25 126.395 ;
			LAYER	M2 ;
			RECT	0 126.295 0.25 126.395 ;
			LAYER	M3 ;
			RECT	0 126.295 0.25 126.395 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[43]

	PIN QA[44]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 129.175 0.25 129.275 ;
			LAYER	M2 ;
			RECT	0 129.175 0.25 129.275 ;
			LAYER	M3 ;
			RECT	0 129.175 0.25 129.275 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[44]

	PIN QA[45]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 132.055 0.25 132.155 ;
			LAYER	M2 ;
			RECT	0 132.055 0.25 132.155 ;
			LAYER	M3 ;
			RECT	0 132.055 0.25 132.155 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[45]

	PIN QA[46]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 134.935 0.25 135.035 ;
			LAYER	M2 ;
			RECT	0 134.935 0.25 135.035 ;
			LAYER	M3 ;
			RECT	0 134.935 0.25 135.035 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[46]

	PIN QA[47]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 137.815 0.25 137.915 ;
			LAYER	M2 ;
			RECT	0 137.815 0.25 137.915 ;
			LAYER	M3 ;
			RECT	0 137.815 0.25 137.915 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[47]

	PIN QA[48]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 140.695 0.25 140.795 ;
			LAYER	M2 ;
			RECT	0 140.695 0.25 140.795 ;
			LAYER	M3 ;
			RECT	0 140.695 0.25 140.795 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[48]

	PIN QA[49]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 143.575 0.25 143.675 ;
			LAYER	M2 ;
			RECT	0 143.575 0.25 143.675 ;
			LAYER	M3 ;
			RECT	0 143.575 0.25 143.675 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[49]

	PIN QA[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 13.975 0.25 14.075 ;
			LAYER	M2 ;
			RECT	0 13.975 0.25 14.075 ;
			LAYER	M3 ;
			RECT	0 13.975 0.25 14.075 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[4]

	PIN QA[50]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 146.455 0.25 146.555 ;
			LAYER	M2 ;
			RECT	0 146.455 0.25 146.555 ;
			LAYER	M3 ;
			RECT	0 146.455 0.25 146.555 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[50]

	PIN QA[51]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 149.335 0.25 149.435 ;
			LAYER	M2 ;
			RECT	0 149.335 0.25 149.435 ;
			LAYER	M3 ;
			RECT	0 149.335 0.25 149.435 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[51]

	PIN QA[52]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 152.215 0.25 152.315 ;
			LAYER	M2 ;
			RECT	0 152.215 0.25 152.315 ;
			LAYER	M3 ;
			RECT	0 152.215 0.25 152.315 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[52]

	PIN QA[53]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 155.095 0.25 155.195 ;
			LAYER	M2 ;
			RECT	0 155.095 0.25 155.195 ;
			LAYER	M3 ;
			RECT	0 155.095 0.25 155.195 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[53]

	PIN QA[54]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 157.975 0.25 158.075 ;
			LAYER	M2 ;
			RECT	0 157.975 0.25 158.075 ;
			LAYER	M3 ;
			RECT	0 157.975 0.25 158.075 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[54]

	PIN QA[55]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 160.855 0.25 160.955 ;
			LAYER	M2 ;
			RECT	0 160.855 0.25 160.955 ;
			LAYER	M3 ;
			RECT	0 160.855 0.25 160.955 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[55]

	PIN QA[56]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 163.735 0.25 163.835 ;
			LAYER	M2 ;
			RECT	0 163.735 0.25 163.835 ;
			LAYER	M3 ;
			RECT	0 163.735 0.25 163.835 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[56]

	PIN QA[57]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 166.615 0.25 166.715 ;
			LAYER	M2 ;
			RECT	0 166.615 0.25 166.715 ;
			LAYER	M3 ;
			RECT	0 166.615 0.25 166.715 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[57]

	PIN QA[58]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 169.495 0.25 169.595 ;
			LAYER	M2 ;
			RECT	0 169.495 0.25 169.595 ;
			LAYER	M3 ;
			RECT	0 169.495 0.25 169.595 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[58]

	PIN QA[59]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 172.375 0.25 172.475 ;
			LAYER	M2 ;
			RECT	0 172.375 0.25 172.475 ;
			LAYER	M3 ;
			RECT	0 172.375 0.25 172.475 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[59]

	PIN QA[5]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 16.855 0.25 16.955 ;
			LAYER	M2 ;
			RECT	0 16.855 0.25 16.955 ;
			LAYER	M3 ;
			RECT	0 16.855 0.25 16.955 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[5]

	PIN QA[60]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 175.255 0.25 175.355 ;
			LAYER	M2 ;
			RECT	0 175.255 0.25 175.355 ;
			LAYER	M3 ;
			RECT	0 175.255 0.25 175.355 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[60]

	PIN QA[61]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 178.135 0.25 178.235 ;
			LAYER	M2 ;
			RECT	0 178.135 0.25 178.235 ;
			LAYER	M3 ;
			RECT	0 178.135 0.25 178.235 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[61]

	PIN QA[62]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 181.015 0.25 181.115 ;
			LAYER	M2 ;
			RECT	0 181.015 0.25 181.115 ;
			LAYER	M3 ;
			RECT	0 181.015 0.25 181.115 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[62]

	PIN QA[63]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 183.895 0.25 183.995 ;
			LAYER	M2 ;
			RECT	0 183.895 0.25 183.995 ;
			LAYER	M3 ;
			RECT	0 183.895 0.25 183.995 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[63]

	PIN QA[64]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 230.865 0.25 230.965 ;
			LAYER	M2 ;
			RECT	0 230.865 0.25 230.965 ;
			LAYER	M3 ;
			RECT	0 230.865 0.25 230.965 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[64]

	PIN QA[65]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 233.745 0.25 233.845 ;
			LAYER	M2 ;
			RECT	0 233.745 0.25 233.845 ;
			LAYER	M3 ;
			RECT	0 233.745 0.25 233.845 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[65]

	PIN QA[66]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 236.625 0.25 236.725 ;
			LAYER	M2 ;
			RECT	0 236.625 0.25 236.725 ;
			LAYER	M3 ;
			RECT	0 236.625 0.25 236.725 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[66]

	PIN QA[67]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 239.505 0.25 239.605 ;
			LAYER	M2 ;
			RECT	0 239.505 0.25 239.605 ;
			LAYER	M3 ;
			RECT	0 239.505 0.25 239.605 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[67]

	PIN QA[68]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 242.385 0.25 242.485 ;
			LAYER	M2 ;
			RECT	0 242.385 0.25 242.485 ;
			LAYER	M3 ;
			RECT	0 242.385 0.25 242.485 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[68]

	PIN QA[69]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 245.265 0.25 245.365 ;
			LAYER	M2 ;
			RECT	0 245.265 0.25 245.365 ;
			LAYER	M3 ;
			RECT	0 245.265 0.25 245.365 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[69]

	PIN QA[6]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 19.735 0.25 19.835 ;
			LAYER	M2 ;
			RECT	0 19.735 0.25 19.835 ;
			LAYER	M3 ;
			RECT	0 19.735 0.25 19.835 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[6]

	PIN QA[70]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 248.145 0.25 248.245 ;
			LAYER	M2 ;
			RECT	0 248.145 0.25 248.245 ;
			LAYER	M3 ;
			RECT	0 248.145 0.25 248.245 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[70]

	PIN QA[71]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 251.025 0.25 251.125 ;
			LAYER	M2 ;
			RECT	0 251.025 0.25 251.125 ;
			LAYER	M3 ;
			RECT	0 251.025 0.25 251.125 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[71]

	PIN QA[72]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 253.905 0.25 254.005 ;
			LAYER	M2 ;
			RECT	0 253.905 0.25 254.005 ;
			LAYER	M3 ;
			RECT	0 253.905 0.25 254.005 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[72]

	PIN QA[73]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 256.785 0.25 256.885 ;
			LAYER	M2 ;
			RECT	0 256.785 0.25 256.885 ;
			LAYER	M3 ;
			RECT	0 256.785 0.25 256.885 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[73]

	PIN QA[74]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 259.665 0.25 259.765 ;
			LAYER	M2 ;
			RECT	0 259.665 0.25 259.765 ;
			LAYER	M3 ;
			RECT	0 259.665 0.25 259.765 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[74]

	PIN QA[75]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 262.545 0.25 262.645 ;
			LAYER	M2 ;
			RECT	0 262.545 0.25 262.645 ;
			LAYER	M3 ;
			RECT	0 262.545 0.25 262.645 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[75]

	PIN QA[76]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 265.425 0.25 265.525 ;
			LAYER	M2 ;
			RECT	0 265.425 0.25 265.525 ;
			LAYER	M3 ;
			RECT	0 265.425 0.25 265.525 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[76]

	PIN QA[77]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 268.305 0.25 268.405 ;
			LAYER	M2 ;
			RECT	0 268.305 0.25 268.405 ;
			LAYER	M3 ;
			RECT	0 268.305 0.25 268.405 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[77]

	PIN QA[78]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 271.185 0.25 271.285 ;
			LAYER	M2 ;
			RECT	0 271.185 0.25 271.285 ;
			LAYER	M3 ;
			RECT	0 271.185 0.25 271.285 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[78]

	PIN QA[79]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 274.065 0.25 274.165 ;
			LAYER	M2 ;
			RECT	0 274.065 0.25 274.165 ;
			LAYER	M3 ;
			RECT	0 274.065 0.25 274.165 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[79]

	PIN QA[7]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 22.615 0.25 22.715 ;
			LAYER	M2 ;
			RECT	0 22.615 0.25 22.715 ;
			LAYER	M3 ;
			RECT	0 22.615 0.25 22.715 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[7]

	PIN QA[80]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 276.945 0.25 277.045 ;
			LAYER	M2 ;
			RECT	0 276.945 0.25 277.045 ;
			LAYER	M3 ;
			RECT	0 276.945 0.25 277.045 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[80]

	PIN QA[81]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 279.825 0.25 279.925 ;
			LAYER	M2 ;
			RECT	0 279.825 0.25 279.925 ;
			LAYER	M3 ;
			RECT	0 279.825 0.25 279.925 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[81]

	PIN QA[82]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 282.705 0.25 282.805 ;
			LAYER	M2 ;
			RECT	0 282.705 0.25 282.805 ;
			LAYER	M3 ;
			RECT	0 282.705 0.25 282.805 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[82]

	PIN QA[83]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 285.585 0.25 285.685 ;
			LAYER	M2 ;
			RECT	0 285.585 0.25 285.685 ;
			LAYER	M3 ;
			RECT	0 285.585 0.25 285.685 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[83]

	PIN QA[84]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 288.465 0.25 288.565 ;
			LAYER	M2 ;
			RECT	0 288.465 0.25 288.565 ;
			LAYER	M3 ;
			RECT	0 288.465 0.25 288.565 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[84]

	PIN QA[85]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 291.345 0.25 291.445 ;
			LAYER	M2 ;
			RECT	0 291.345 0.25 291.445 ;
			LAYER	M3 ;
			RECT	0 291.345 0.25 291.445 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[85]

	PIN QA[86]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 294.225 0.25 294.325 ;
			LAYER	M2 ;
			RECT	0 294.225 0.25 294.325 ;
			LAYER	M3 ;
			RECT	0 294.225 0.25 294.325 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[86]

	PIN QA[87]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 297.105 0.25 297.205 ;
			LAYER	M2 ;
			RECT	0 297.105 0.25 297.205 ;
			LAYER	M3 ;
			RECT	0 297.105 0.25 297.205 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[87]

	PIN QA[88]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 299.985 0.25 300.085 ;
			LAYER	M2 ;
			RECT	0 299.985 0.25 300.085 ;
			LAYER	M3 ;
			RECT	0 299.985 0.25 300.085 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[88]

	PIN QA[89]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 302.865 0.25 302.965 ;
			LAYER	M2 ;
			RECT	0 302.865 0.25 302.965 ;
			LAYER	M3 ;
			RECT	0 302.865 0.25 302.965 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[89]

	PIN QA[8]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 25.495 0.25 25.595 ;
			LAYER	M2 ;
			RECT	0 25.495 0.25 25.595 ;
			LAYER	M3 ;
			RECT	0 25.495 0.25 25.595 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[8]

	PIN QA[90]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 305.745 0.25 305.845 ;
			LAYER	M2 ;
			RECT	0 305.745 0.25 305.845 ;
			LAYER	M3 ;
			RECT	0 305.745 0.25 305.845 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[90]

	PIN QA[91]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 308.625 0.25 308.725 ;
			LAYER	M2 ;
			RECT	0 308.625 0.25 308.725 ;
			LAYER	M3 ;
			RECT	0 308.625 0.25 308.725 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[91]

	PIN QA[92]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 311.505 0.25 311.605 ;
			LAYER	M2 ;
			RECT	0 311.505 0.25 311.605 ;
			LAYER	M3 ;
			RECT	0 311.505 0.25 311.605 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[92]

	PIN QA[93]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 314.385 0.25 314.485 ;
			LAYER	M2 ;
			RECT	0 314.385 0.25 314.485 ;
			LAYER	M3 ;
			RECT	0 314.385 0.25 314.485 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[93]

	PIN QA[94]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 317.265 0.25 317.365 ;
			LAYER	M2 ;
			RECT	0 317.265 0.25 317.365 ;
			LAYER	M3 ;
			RECT	0 317.265 0.25 317.365 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[94]

	PIN QA[95]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 320.145 0.25 320.245 ;
			LAYER	M2 ;
			RECT	0 320.145 0.25 320.245 ;
			LAYER	M3 ;
			RECT	0 320.145 0.25 320.245 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[95]

	PIN QA[96]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 323.025 0.25 323.125 ;
			LAYER	M2 ;
			RECT	0 323.025 0.25 323.125 ;
			LAYER	M3 ;
			RECT	0 323.025 0.25 323.125 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[96]

	PIN QA[97]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 325.905 0.25 326.005 ;
			LAYER	M2 ;
			RECT	0 325.905 0.25 326.005 ;
			LAYER	M3 ;
			RECT	0 325.905 0.25 326.005 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[97]

	PIN QA[98]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 328.785 0.25 328.885 ;
			LAYER	M2 ;
			RECT	0 328.785 0.25 328.885 ;
			LAYER	M3 ;
			RECT	0 328.785 0.25 328.885 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[98]

	PIN QA[99]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 331.665 0.25 331.765 ;
			LAYER	M2 ;
			RECT	0 331.665 0.25 331.765 ;
			LAYER	M3 ;
			RECT	0 331.665 0.25 331.765 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[99]

	PIN QA[9]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 28.375 0.25 28.475 ;
			LAYER	M2 ;
			RECT	0 28.375 0.25 28.475 ;
			LAYER	M3 ;
			RECT	0 28.375 0.25 28.475 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[9]

	PIN RET1N
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 188.11 0.25 188.21 ;
			LAYER	M2 ;
			RECT	0 188.11 0.25 188.21 ;
			LAYER	M3 ;
			RECT	0 188.11 0.25 188.21 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END RET1N

	PIN SEA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 205.9 0.25 206 ;
			LAYER	M2 ;
			RECT	0 205.9 0.25 206 ;
			LAYER	M3 ;
			RECT	0 205.9 0.25 206 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SEA

	PIN SEB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 208.735 0.25 208.835 ;
			LAYER	M2 ;
			RECT	0 208.735 0.25 208.835 ;
			LAYER	M3 ;
			RECT	0 208.735 0.25 208.835 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SEB

	PIN SIA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 206.1 0.25 206.2 ;
			LAYER	M2 ;
			RECT	0 206.1 0.25 206.2 ;
			LAYER	M3 ;
			RECT	0 206.1 0.25 206.2 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIA[0]

	PIN SIA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 207.07 0.25 207.17 ;
			LAYER	M2 ;
			RECT	0 207.07 0.25 207.17 ;
			LAYER	M3 ;
			RECT	0 207.07 0.25 207.17 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIA[1]

	PIN SIB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 202.675 0.25 202.775 ;
			LAYER	M2 ;
			RECT	0 202.675 0.25 202.775 ;
			LAYER	M3 ;
			RECT	0 202.675 0.25 202.775 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIB[0]

	PIN SIB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 220.325 0.25 220.425 ;
			LAYER	M2 ;
			RECT	0 220.325 0.25 220.425 ;
			LAYER	M3 ;
			RECT	0 220.325 0.25 220.425 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIB[1]

	PIN SOA[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 0.36 0.25 0.46 ;
			LAYER	M2 ;
			RECT	0 0.36 0.25 0.46 ;
			LAYER	M3 ;
			RECT	0 0.36 0.25 0.46 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOA[0]

	PIN SOA[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 414.4 0.25 414.5 ;
			LAYER	M2 ;
			RECT	0 414.4 0.25 414.5 ;
			LAYER	M3 ;
			RECT	0 414.4 0.25 414.5 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOA[1]

	PIN SOB[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 0.09 0.25 0.19 ;
			LAYER	M2 ;
			RECT	0 0.09 0.25 0.19 ;
			LAYER	M3 ;
			RECT	0 0.09 0.25 0.19 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOB[0]

	PIN SOB[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 414.67 0.25 414.77 ;
			LAYER	M2 ;
			RECT	0 414.67 0.25 414.77 ;
			LAYER	M3 ;
			RECT	0 414.67 0.25 414.77 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOB[1]

	PIN TAA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 190.755 0.25 190.855 ;
			LAYER	M2 ;
			RECT	0 190.755 0.25 190.855 ;
			LAYER	M3 ;
			RECT	0 190.755 0.25 190.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[0]

	PIN TAA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 193.785 0.25 193.885 ;
			LAYER	M2 ;
			RECT	0 193.785 0.25 193.885 ;
			LAYER	M3 ;
			RECT	0 193.785 0.25 193.885 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[1]

	PIN TAA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 196.845 0.25 196.945 ;
			LAYER	M2 ;
			RECT	0 196.845 0.25 196.945 ;
			LAYER	M3 ;
			RECT	0 196.845 0.25 196.945 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[2]

	PIN TAA[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 199.36 0.25 199.46 ;
			LAYER	M2 ;
			RECT	0 199.36 0.25 199.46 ;
			LAYER	M3 ;
			RECT	0 199.36 0.25 199.46 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[3]

	PIN TAA[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 202.39 0.25 202.49 ;
			LAYER	M2 ;
			RECT	0 202.39 0.25 202.49 ;
			LAYER	M3 ;
			RECT	0 202.39 0.25 202.49 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[4]

	PIN TAB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 224.67 0.25 224.77 ;
			LAYER	M2 ;
			RECT	0 224.67 0.25 224.77 ;
			LAYER	M3 ;
			RECT	0 224.67 0.25 224.77 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[0]

	PIN TAB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 221.64 0.25 221.74 ;
			LAYER	M2 ;
			RECT	0 221.64 0.25 221.74 ;
			LAYER	M3 ;
			RECT	0 221.64 0.25 221.74 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[1]

	PIN TAB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 218.58 0.25 218.68 ;
			LAYER	M2 ;
			RECT	0 218.58 0.25 218.68 ;
			LAYER	M3 ;
			RECT	0 218.58 0.25 218.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[2]

	PIN TAB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 216.095 0.25 216.195 ;
			LAYER	M2 ;
			RECT	0 216.095 0.25 216.195 ;
			LAYER	M3 ;
			RECT	0 216.095 0.25 216.195 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[3]

	PIN TAB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 213.06 0.25 213.16 ;
			LAYER	M2 ;
			RECT	0 213.06 0.25 213.16 ;
			LAYER	M3 ;
			RECT	0 213.06 0.25 213.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[4]

	PIN TCENA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 188.31 0.25 188.41 ;
			LAYER	M2 ;
			RECT	0 188.31 0.25 188.41 ;
			LAYER	M3 ;
			RECT	0 188.31 0.25 188.41 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TCENA

	PIN TCENB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 228.31 0.25 228.41 ;
			LAYER	M2 ;
			RECT	0 228.31 0.25 228.41 ;
			LAYER	M3 ;
			RECT	0 228.31 0.25 228.41 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TCENB

	PIN TDB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 1.465 0.25 1.565 ;
			LAYER	M2 ;
			RECT	0 1.465 0.25 1.565 ;
			LAYER	M3 ;
			RECT	0 1.465 0.25 1.565 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[0]

	PIN TDB[100]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 335.535 0.25 335.635 ;
			LAYER	M2 ;
			RECT	0 335.535 0.25 335.635 ;
			LAYER	M3 ;
			RECT	0 335.535 0.25 335.635 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[100]

	PIN TDB[101]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 338.415 0.25 338.515 ;
			LAYER	M2 ;
			RECT	0 338.415 0.25 338.515 ;
			LAYER	M3 ;
			RECT	0 338.415 0.25 338.515 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[101]

	PIN TDB[102]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 341.295 0.25 341.395 ;
			LAYER	M2 ;
			RECT	0 341.295 0.25 341.395 ;
			LAYER	M3 ;
			RECT	0 341.295 0.25 341.395 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[102]

	PIN TDB[103]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 344.175 0.25 344.275 ;
			LAYER	M2 ;
			RECT	0 344.175 0.25 344.275 ;
			LAYER	M3 ;
			RECT	0 344.175 0.25 344.275 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[103]

	PIN TDB[104]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 347.055 0.25 347.155 ;
			LAYER	M2 ;
			RECT	0 347.055 0.25 347.155 ;
			LAYER	M3 ;
			RECT	0 347.055 0.25 347.155 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[104]

	PIN TDB[105]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 349.935 0.25 350.035 ;
			LAYER	M2 ;
			RECT	0 349.935 0.25 350.035 ;
			LAYER	M3 ;
			RECT	0 349.935 0.25 350.035 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[105]

	PIN TDB[106]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 352.815 0.25 352.915 ;
			LAYER	M2 ;
			RECT	0 352.815 0.25 352.915 ;
			LAYER	M3 ;
			RECT	0 352.815 0.25 352.915 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[106]

	PIN TDB[107]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 355.695 0.25 355.795 ;
			LAYER	M2 ;
			RECT	0 355.695 0.25 355.795 ;
			LAYER	M3 ;
			RECT	0 355.695 0.25 355.795 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[107]

	PIN TDB[108]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 358.575 0.25 358.675 ;
			LAYER	M2 ;
			RECT	0 358.575 0.25 358.675 ;
			LAYER	M3 ;
			RECT	0 358.575 0.25 358.675 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[108]

	PIN TDB[109]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 361.455 0.25 361.555 ;
			LAYER	M2 ;
			RECT	0 361.455 0.25 361.555 ;
			LAYER	M3 ;
			RECT	0 361.455 0.25 361.555 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[109]

	PIN TDB[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 30.265 0.25 30.365 ;
			LAYER	M2 ;
			RECT	0 30.265 0.25 30.365 ;
			LAYER	M3 ;
			RECT	0 30.265 0.25 30.365 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[10]

	PIN TDB[110]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 364.335 0.25 364.435 ;
			LAYER	M2 ;
			RECT	0 364.335 0.25 364.435 ;
			LAYER	M3 ;
			RECT	0 364.335 0.25 364.435 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[110]

	PIN TDB[111]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 367.215 0.25 367.315 ;
			LAYER	M2 ;
			RECT	0 367.215 0.25 367.315 ;
			LAYER	M3 ;
			RECT	0 367.215 0.25 367.315 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[111]

	PIN TDB[112]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 370.095 0.25 370.195 ;
			LAYER	M2 ;
			RECT	0 370.095 0.25 370.195 ;
			LAYER	M3 ;
			RECT	0 370.095 0.25 370.195 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[112]

	PIN TDB[113]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 372.975 0.25 373.075 ;
			LAYER	M2 ;
			RECT	0 372.975 0.25 373.075 ;
			LAYER	M3 ;
			RECT	0 372.975 0.25 373.075 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[113]

	PIN TDB[114]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 375.855 0.25 375.955 ;
			LAYER	M2 ;
			RECT	0 375.855 0.25 375.955 ;
			LAYER	M3 ;
			RECT	0 375.855 0.25 375.955 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[114]

	PIN TDB[115]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 378.735 0.25 378.835 ;
			LAYER	M2 ;
			RECT	0 378.735 0.25 378.835 ;
			LAYER	M3 ;
			RECT	0 378.735 0.25 378.835 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[115]

	PIN TDB[116]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 381.615 0.25 381.715 ;
			LAYER	M2 ;
			RECT	0 381.615 0.25 381.715 ;
			LAYER	M3 ;
			RECT	0 381.615 0.25 381.715 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[116]

	PIN TDB[117]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 384.495 0.25 384.595 ;
			LAYER	M2 ;
			RECT	0 384.495 0.25 384.595 ;
			LAYER	M3 ;
			RECT	0 384.495 0.25 384.595 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[117]

	PIN TDB[118]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 387.375 0.25 387.475 ;
			LAYER	M2 ;
			RECT	0 387.375 0.25 387.475 ;
			LAYER	M3 ;
			RECT	0 387.375 0.25 387.475 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[118]

	PIN TDB[119]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 390.255 0.25 390.355 ;
			LAYER	M2 ;
			RECT	0 390.255 0.25 390.355 ;
			LAYER	M3 ;
			RECT	0 390.255 0.25 390.355 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[119]

	PIN TDB[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 33.145 0.25 33.245 ;
			LAYER	M2 ;
			RECT	0 33.145 0.25 33.245 ;
			LAYER	M3 ;
			RECT	0 33.145 0.25 33.245 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[11]

	PIN TDB[120]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 393.135 0.25 393.235 ;
			LAYER	M2 ;
			RECT	0 393.135 0.25 393.235 ;
			LAYER	M3 ;
			RECT	0 393.135 0.25 393.235 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[120]

	PIN TDB[121]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 396.015 0.25 396.115 ;
			LAYER	M2 ;
			RECT	0 396.015 0.25 396.115 ;
			LAYER	M3 ;
			RECT	0 396.015 0.25 396.115 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[121]

	PIN TDB[122]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 398.895 0.25 398.995 ;
			LAYER	M2 ;
			RECT	0 398.895 0.25 398.995 ;
			LAYER	M3 ;
			RECT	0 398.895 0.25 398.995 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[122]

	PIN TDB[123]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 401.775 0.25 401.875 ;
			LAYER	M2 ;
			RECT	0 401.775 0.25 401.875 ;
			LAYER	M3 ;
			RECT	0 401.775 0.25 401.875 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[123]

	PIN TDB[124]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 404.655 0.25 404.755 ;
			LAYER	M2 ;
			RECT	0 404.655 0.25 404.755 ;
			LAYER	M3 ;
			RECT	0 404.655 0.25 404.755 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[124]

	PIN TDB[125]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 407.535 0.25 407.635 ;
			LAYER	M2 ;
			RECT	0 407.535 0.25 407.635 ;
			LAYER	M3 ;
			RECT	0 407.535 0.25 407.635 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[125]

	PIN TDB[126]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 410.415 0.25 410.515 ;
			LAYER	M2 ;
			RECT	0 410.415 0.25 410.515 ;
			LAYER	M3 ;
			RECT	0 410.415 0.25 410.515 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[126]

	PIN TDB[127]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 413.295 0.25 413.395 ;
			LAYER	M2 ;
			RECT	0 413.295 0.25 413.395 ;
			LAYER	M3 ;
			RECT	0 413.295 0.25 413.395 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[127]

	PIN TDB[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 36.025 0.25 36.125 ;
			LAYER	M2 ;
			RECT	0 36.025 0.25 36.125 ;
			LAYER	M3 ;
			RECT	0 36.025 0.25 36.125 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[12]

	PIN TDB[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 38.905 0.25 39.005 ;
			LAYER	M2 ;
			RECT	0 38.905 0.25 39.005 ;
			LAYER	M3 ;
			RECT	0 38.905 0.25 39.005 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[13]

	PIN TDB[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 41.785 0.25 41.885 ;
			LAYER	M2 ;
			RECT	0 41.785 0.25 41.885 ;
			LAYER	M3 ;
			RECT	0 41.785 0.25 41.885 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[14]

	PIN TDB[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 44.665 0.25 44.765 ;
			LAYER	M2 ;
			RECT	0 44.665 0.25 44.765 ;
			LAYER	M3 ;
			RECT	0 44.665 0.25 44.765 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[15]

	PIN TDB[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 47.545 0.25 47.645 ;
			LAYER	M2 ;
			RECT	0 47.545 0.25 47.645 ;
			LAYER	M3 ;
			RECT	0 47.545 0.25 47.645 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[16]

	PIN TDB[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 50.425 0.25 50.525 ;
			LAYER	M2 ;
			RECT	0 50.425 0.25 50.525 ;
			LAYER	M3 ;
			RECT	0 50.425 0.25 50.525 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[17]

	PIN TDB[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 53.305 0.25 53.405 ;
			LAYER	M2 ;
			RECT	0 53.305 0.25 53.405 ;
			LAYER	M3 ;
			RECT	0 53.305 0.25 53.405 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[18]

	PIN TDB[19]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 56.185 0.25 56.285 ;
			LAYER	M2 ;
			RECT	0 56.185 0.25 56.285 ;
			LAYER	M3 ;
			RECT	0 56.185 0.25 56.285 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[19]

	PIN TDB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 4.345 0.25 4.445 ;
			LAYER	M2 ;
			RECT	0 4.345 0.25 4.445 ;
			LAYER	M3 ;
			RECT	0 4.345 0.25 4.445 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[1]

	PIN TDB[20]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 59.065 0.25 59.165 ;
			LAYER	M2 ;
			RECT	0 59.065 0.25 59.165 ;
			LAYER	M3 ;
			RECT	0 59.065 0.25 59.165 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[20]

	PIN TDB[21]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 61.945 0.25 62.045 ;
			LAYER	M2 ;
			RECT	0 61.945 0.25 62.045 ;
			LAYER	M3 ;
			RECT	0 61.945 0.25 62.045 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[21]

	PIN TDB[22]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 64.825 0.25 64.925 ;
			LAYER	M2 ;
			RECT	0 64.825 0.25 64.925 ;
			LAYER	M3 ;
			RECT	0 64.825 0.25 64.925 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[22]

	PIN TDB[23]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 67.705 0.25 67.805 ;
			LAYER	M2 ;
			RECT	0 67.705 0.25 67.805 ;
			LAYER	M3 ;
			RECT	0 67.705 0.25 67.805 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[23]

	PIN TDB[24]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 70.585 0.25 70.685 ;
			LAYER	M2 ;
			RECT	0 70.585 0.25 70.685 ;
			LAYER	M3 ;
			RECT	0 70.585 0.25 70.685 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[24]

	PIN TDB[25]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 73.465 0.25 73.565 ;
			LAYER	M2 ;
			RECT	0 73.465 0.25 73.565 ;
			LAYER	M3 ;
			RECT	0 73.465 0.25 73.565 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[25]

	PIN TDB[26]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 76.345 0.25 76.445 ;
			LAYER	M2 ;
			RECT	0 76.345 0.25 76.445 ;
			LAYER	M3 ;
			RECT	0 76.345 0.25 76.445 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[26]

	PIN TDB[27]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 79.225 0.25 79.325 ;
			LAYER	M2 ;
			RECT	0 79.225 0.25 79.325 ;
			LAYER	M3 ;
			RECT	0 79.225 0.25 79.325 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[27]

	PIN TDB[28]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 82.105 0.25 82.205 ;
			LAYER	M2 ;
			RECT	0 82.105 0.25 82.205 ;
			LAYER	M3 ;
			RECT	0 82.105 0.25 82.205 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[28]

	PIN TDB[29]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 84.985 0.25 85.085 ;
			LAYER	M2 ;
			RECT	0 84.985 0.25 85.085 ;
			LAYER	M3 ;
			RECT	0 84.985 0.25 85.085 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[29]

	PIN TDB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 7.225 0.25 7.325 ;
			LAYER	M2 ;
			RECT	0 7.225 0.25 7.325 ;
			LAYER	M3 ;
			RECT	0 7.225 0.25 7.325 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[2]

	PIN TDB[30]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 87.865 0.25 87.965 ;
			LAYER	M2 ;
			RECT	0 87.865 0.25 87.965 ;
			LAYER	M3 ;
			RECT	0 87.865 0.25 87.965 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[30]

	PIN TDB[31]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 90.745 0.25 90.845 ;
			LAYER	M2 ;
			RECT	0 90.745 0.25 90.845 ;
			LAYER	M3 ;
			RECT	0 90.745 0.25 90.845 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[31]

	PIN TDB[32]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 93.625 0.25 93.725 ;
			LAYER	M2 ;
			RECT	0 93.625 0.25 93.725 ;
			LAYER	M3 ;
			RECT	0 93.625 0.25 93.725 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[32]

	PIN TDB[33]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 96.505 0.25 96.605 ;
			LAYER	M2 ;
			RECT	0 96.505 0.25 96.605 ;
			LAYER	M3 ;
			RECT	0 96.505 0.25 96.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[33]

	PIN TDB[34]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 99.385 0.25 99.485 ;
			LAYER	M2 ;
			RECT	0 99.385 0.25 99.485 ;
			LAYER	M3 ;
			RECT	0 99.385 0.25 99.485 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[34]

	PIN TDB[35]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 102.265 0.25 102.365 ;
			LAYER	M2 ;
			RECT	0 102.265 0.25 102.365 ;
			LAYER	M3 ;
			RECT	0 102.265 0.25 102.365 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[35]

	PIN TDB[36]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 105.145 0.25 105.245 ;
			LAYER	M2 ;
			RECT	0 105.145 0.25 105.245 ;
			LAYER	M3 ;
			RECT	0 105.145 0.25 105.245 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[36]

	PIN TDB[37]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 108.025 0.25 108.125 ;
			LAYER	M2 ;
			RECT	0 108.025 0.25 108.125 ;
			LAYER	M3 ;
			RECT	0 108.025 0.25 108.125 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[37]

	PIN TDB[38]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 110.905 0.25 111.005 ;
			LAYER	M2 ;
			RECT	0 110.905 0.25 111.005 ;
			LAYER	M3 ;
			RECT	0 110.905 0.25 111.005 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[38]

	PIN TDB[39]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 113.785 0.25 113.885 ;
			LAYER	M2 ;
			RECT	0 113.785 0.25 113.885 ;
			LAYER	M3 ;
			RECT	0 113.785 0.25 113.885 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[39]

	PIN TDB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 10.105 0.25 10.205 ;
			LAYER	M2 ;
			RECT	0 10.105 0.25 10.205 ;
			LAYER	M3 ;
			RECT	0 10.105 0.25 10.205 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[3]

	PIN TDB[40]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 116.665 0.25 116.765 ;
			LAYER	M2 ;
			RECT	0 116.665 0.25 116.765 ;
			LAYER	M3 ;
			RECT	0 116.665 0.25 116.765 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[40]

	PIN TDB[41]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 119.545 0.25 119.645 ;
			LAYER	M2 ;
			RECT	0 119.545 0.25 119.645 ;
			LAYER	M3 ;
			RECT	0 119.545 0.25 119.645 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[41]

	PIN TDB[42]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 122.425 0.25 122.525 ;
			LAYER	M2 ;
			RECT	0 122.425 0.25 122.525 ;
			LAYER	M3 ;
			RECT	0 122.425 0.25 122.525 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[42]

	PIN TDB[43]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 125.305 0.25 125.405 ;
			LAYER	M2 ;
			RECT	0 125.305 0.25 125.405 ;
			LAYER	M3 ;
			RECT	0 125.305 0.25 125.405 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[43]

	PIN TDB[44]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 128.185 0.25 128.285 ;
			LAYER	M2 ;
			RECT	0 128.185 0.25 128.285 ;
			LAYER	M3 ;
			RECT	0 128.185 0.25 128.285 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[44]

	PIN TDB[45]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 131.065 0.25 131.165 ;
			LAYER	M2 ;
			RECT	0 131.065 0.25 131.165 ;
			LAYER	M3 ;
			RECT	0 131.065 0.25 131.165 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[45]

	PIN TDB[46]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 133.945 0.25 134.045 ;
			LAYER	M2 ;
			RECT	0 133.945 0.25 134.045 ;
			LAYER	M3 ;
			RECT	0 133.945 0.25 134.045 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[46]

	PIN TDB[47]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 136.825 0.25 136.925 ;
			LAYER	M2 ;
			RECT	0 136.825 0.25 136.925 ;
			LAYER	M3 ;
			RECT	0 136.825 0.25 136.925 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[47]

	PIN TDB[48]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 139.705 0.25 139.805 ;
			LAYER	M2 ;
			RECT	0 139.705 0.25 139.805 ;
			LAYER	M3 ;
			RECT	0 139.705 0.25 139.805 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[48]

	PIN TDB[49]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 142.585 0.25 142.685 ;
			LAYER	M2 ;
			RECT	0 142.585 0.25 142.685 ;
			LAYER	M3 ;
			RECT	0 142.585 0.25 142.685 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[49]

	PIN TDB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 12.985 0.25 13.085 ;
			LAYER	M2 ;
			RECT	0 12.985 0.25 13.085 ;
			LAYER	M3 ;
			RECT	0 12.985 0.25 13.085 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[4]

	PIN TDB[50]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 145.465 0.25 145.565 ;
			LAYER	M2 ;
			RECT	0 145.465 0.25 145.565 ;
			LAYER	M3 ;
			RECT	0 145.465 0.25 145.565 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[50]

	PIN TDB[51]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 148.345 0.25 148.445 ;
			LAYER	M2 ;
			RECT	0 148.345 0.25 148.445 ;
			LAYER	M3 ;
			RECT	0 148.345 0.25 148.445 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[51]

	PIN TDB[52]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 151.225 0.25 151.325 ;
			LAYER	M2 ;
			RECT	0 151.225 0.25 151.325 ;
			LAYER	M3 ;
			RECT	0 151.225 0.25 151.325 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[52]

	PIN TDB[53]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 154.105 0.25 154.205 ;
			LAYER	M2 ;
			RECT	0 154.105 0.25 154.205 ;
			LAYER	M3 ;
			RECT	0 154.105 0.25 154.205 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[53]

	PIN TDB[54]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 156.985 0.25 157.085 ;
			LAYER	M2 ;
			RECT	0 156.985 0.25 157.085 ;
			LAYER	M3 ;
			RECT	0 156.985 0.25 157.085 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[54]

	PIN TDB[55]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 159.865 0.25 159.965 ;
			LAYER	M2 ;
			RECT	0 159.865 0.25 159.965 ;
			LAYER	M3 ;
			RECT	0 159.865 0.25 159.965 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[55]

	PIN TDB[56]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 162.745 0.25 162.845 ;
			LAYER	M2 ;
			RECT	0 162.745 0.25 162.845 ;
			LAYER	M3 ;
			RECT	0 162.745 0.25 162.845 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[56]

	PIN TDB[57]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 165.625 0.25 165.725 ;
			LAYER	M2 ;
			RECT	0 165.625 0.25 165.725 ;
			LAYER	M3 ;
			RECT	0 165.625 0.25 165.725 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[57]

	PIN TDB[58]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 168.505 0.25 168.605 ;
			LAYER	M2 ;
			RECT	0 168.505 0.25 168.605 ;
			LAYER	M3 ;
			RECT	0 168.505 0.25 168.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[58]

	PIN TDB[59]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 171.385 0.25 171.485 ;
			LAYER	M2 ;
			RECT	0 171.385 0.25 171.485 ;
			LAYER	M3 ;
			RECT	0 171.385 0.25 171.485 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[59]

	PIN TDB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 15.865 0.25 15.965 ;
			LAYER	M2 ;
			RECT	0 15.865 0.25 15.965 ;
			LAYER	M3 ;
			RECT	0 15.865 0.25 15.965 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[5]

	PIN TDB[60]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 174.265 0.25 174.365 ;
			LAYER	M2 ;
			RECT	0 174.265 0.25 174.365 ;
			LAYER	M3 ;
			RECT	0 174.265 0.25 174.365 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[60]

	PIN TDB[61]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 177.145 0.25 177.245 ;
			LAYER	M2 ;
			RECT	0 177.145 0.25 177.245 ;
			LAYER	M3 ;
			RECT	0 177.145 0.25 177.245 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[61]

	PIN TDB[62]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 180.025 0.25 180.125 ;
			LAYER	M2 ;
			RECT	0 180.025 0.25 180.125 ;
			LAYER	M3 ;
			RECT	0 180.025 0.25 180.125 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[62]

	PIN TDB[63]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 182.905 0.25 183.005 ;
			LAYER	M2 ;
			RECT	0 182.905 0.25 183.005 ;
			LAYER	M3 ;
			RECT	0 182.905 0.25 183.005 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[63]

	PIN TDB[64]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 231.855 0.25 231.955 ;
			LAYER	M2 ;
			RECT	0 231.855 0.25 231.955 ;
			LAYER	M3 ;
			RECT	0 231.855 0.25 231.955 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[64]

	PIN TDB[65]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 234.735 0.25 234.835 ;
			LAYER	M2 ;
			RECT	0 234.735 0.25 234.835 ;
			LAYER	M3 ;
			RECT	0 234.735 0.25 234.835 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[65]

	PIN TDB[66]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 237.615 0.25 237.715 ;
			LAYER	M2 ;
			RECT	0 237.615 0.25 237.715 ;
			LAYER	M3 ;
			RECT	0 237.615 0.25 237.715 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[66]

	PIN TDB[67]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 240.495 0.25 240.595 ;
			LAYER	M2 ;
			RECT	0 240.495 0.25 240.595 ;
			LAYER	M3 ;
			RECT	0 240.495 0.25 240.595 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[67]

	PIN TDB[68]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 243.375 0.25 243.475 ;
			LAYER	M2 ;
			RECT	0 243.375 0.25 243.475 ;
			LAYER	M3 ;
			RECT	0 243.375 0.25 243.475 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[68]

	PIN TDB[69]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 246.255 0.25 246.355 ;
			LAYER	M2 ;
			RECT	0 246.255 0.25 246.355 ;
			LAYER	M3 ;
			RECT	0 246.255 0.25 246.355 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[69]

	PIN TDB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 18.745 0.25 18.845 ;
			LAYER	M2 ;
			RECT	0 18.745 0.25 18.845 ;
			LAYER	M3 ;
			RECT	0 18.745 0.25 18.845 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[6]

	PIN TDB[70]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 249.135 0.25 249.235 ;
			LAYER	M2 ;
			RECT	0 249.135 0.25 249.235 ;
			LAYER	M3 ;
			RECT	0 249.135 0.25 249.235 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[70]

	PIN TDB[71]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 252.015 0.25 252.115 ;
			LAYER	M2 ;
			RECT	0 252.015 0.25 252.115 ;
			LAYER	M3 ;
			RECT	0 252.015 0.25 252.115 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[71]

	PIN TDB[72]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 254.895 0.25 254.995 ;
			LAYER	M2 ;
			RECT	0 254.895 0.25 254.995 ;
			LAYER	M3 ;
			RECT	0 254.895 0.25 254.995 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[72]

	PIN TDB[73]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 257.775 0.25 257.875 ;
			LAYER	M2 ;
			RECT	0 257.775 0.25 257.875 ;
			LAYER	M3 ;
			RECT	0 257.775 0.25 257.875 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[73]

	PIN TDB[74]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 260.655 0.25 260.755 ;
			LAYER	M2 ;
			RECT	0 260.655 0.25 260.755 ;
			LAYER	M3 ;
			RECT	0 260.655 0.25 260.755 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[74]

	PIN TDB[75]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 263.535 0.25 263.635 ;
			LAYER	M2 ;
			RECT	0 263.535 0.25 263.635 ;
			LAYER	M3 ;
			RECT	0 263.535 0.25 263.635 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[75]

	PIN TDB[76]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 266.415 0.25 266.515 ;
			LAYER	M2 ;
			RECT	0 266.415 0.25 266.515 ;
			LAYER	M3 ;
			RECT	0 266.415 0.25 266.515 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[76]

	PIN TDB[77]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 269.295 0.25 269.395 ;
			LAYER	M2 ;
			RECT	0 269.295 0.25 269.395 ;
			LAYER	M3 ;
			RECT	0 269.295 0.25 269.395 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[77]

	PIN TDB[78]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 272.175 0.25 272.275 ;
			LAYER	M2 ;
			RECT	0 272.175 0.25 272.275 ;
			LAYER	M3 ;
			RECT	0 272.175 0.25 272.275 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[78]

	PIN TDB[79]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 275.055 0.25 275.155 ;
			LAYER	M2 ;
			RECT	0 275.055 0.25 275.155 ;
			LAYER	M3 ;
			RECT	0 275.055 0.25 275.155 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[79]

	PIN TDB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 21.625 0.25 21.725 ;
			LAYER	M2 ;
			RECT	0 21.625 0.25 21.725 ;
			LAYER	M3 ;
			RECT	0 21.625 0.25 21.725 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[7]

	PIN TDB[80]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 277.935 0.25 278.035 ;
			LAYER	M2 ;
			RECT	0 277.935 0.25 278.035 ;
			LAYER	M3 ;
			RECT	0 277.935 0.25 278.035 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[80]

	PIN TDB[81]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 280.815 0.25 280.915 ;
			LAYER	M2 ;
			RECT	0 280.815 0.25 280.915 ;
			LAYER	M3 ;
			RECT	0 280.815 0.25 280.915 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[81]

	PIN TDB[82]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 283.695 0.25 283.795 ;
			LAYER	M2 ;
			RECT	0 283.695 0.25 283.795 ;
			LAYER	M3 ;
			RECT	0 283.695 0.25 283.795 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[82]

	PIN TDB[83]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 286.575 0.25 286.675 ;
			LAYER	M2 ;
			RECT	0 286.575 0.25 286.675 ;
			LAYER	M3 ;
			RECT	0 286.575 0.25 286.675 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[83]

	PIN TDB[84]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 289.455 0.25 289.555 ;
			LAYER	M2 ;
			RECT	0 289.455 0.25 289.555 ;
			LAYER	M3 ;
			RECT	0 289.455 0.25 289.555 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[84]

	PIN TDB[85]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 292.335 0.25 292.435 ;
			LAYER	M2 ;
			RECT	0 292.335 0.25 292.435 ;
			LAYER	M3 ;
			RECT	0 292.335 0.25 292.435 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[85]

	PIN TDB[86]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 295.215 0.25 295.315 ;
			LAYER	M2 ;
			RECT	0 295.215 0.25 295.315 ;
			LAYER	M3 ;
			RECT	0 295.215 0.25 295.315 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[86]

	PIN TDB[87]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 298.095 0.25 298.195 ;
			LAYER	M2 ;
			RECT	0 298.095 0.25 298.195 ;
			LAYER	M3 ;
			RECT	0 298.095 0.25 298.195 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[87]

	PIN TDB[88]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 300.975 0.25 301.075 ;
			LAYER	M2 ;
			RECT	0 300.975 0.25 301.075 ;
			LAYER	M3 ;
			RECT	0 300.975 0.25 301.075 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[88]

	PIN TDB[89]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 303.855 0.25 303.955 ;
			LAYER	M2 ;
			RECT	0 303.855 0.25 303.955 ;
			LAYER	M3 ;
			RECT	0 303.855 0.25 303.955 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[89]

	PIN TDB[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 24.505 0.25 24.605 ;
			LAYER	M2 ;
			RECT	0 24.505 0.25 24.605 ;
			LAYER	M3 ;
			RECT	0 24.505 0.25 24.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[8]

	PIN TDB[90]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 306.735 0.25 306.835 ;
			LAYER	M2 ;
			RECT	0 306.735 0.25 306.835 ;
			LAYER	M3 ;
			RECT	0 306.735 0.25 306.835 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[90]

	PIN TDB[91]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 309.615 0.25 309.715 ;
			LAYER	M2 ;
			RECT	0 309.615 0.25 309.715 ;
			LAYER	M3 ;
			RECT	0 309.615 0.25 309.715 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[91]

	PIN TDB[92]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 312.495 0.25 312.595 ;
			LAYER	M2 ;
			RECT	0 312.495 0.25 312.595 ;
			LAYER	M3 ;
			RECT	0 312.495 0.25 312.595 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[92]

	PIN TDB[93]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 315.375 0.25 315.475 ;
			LAYER	M2 ;
			RECT	0 315.375 0.25 315.475 ;
			LAYER	M3 ;
			RECT	0 315.375 0.25 315.475 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[93]

	PIN TDB[94]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 318.255 0.25 318.355 ;
			LAYER	M2 ;
			RECT	0 318.255 0.25 318.355 ;
			LAYER	M3 ;
			RECT	0 318.255 0.25 318.355 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[94]

	PIN TDB[95]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 321.135 0.25 321.235 ;
			LAYER	M2 ;
			RECT	0 321.135 0.25 321.235 ;
			LAYER	M3 ;
			RECT	0 321.135 0.25 321.235 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[95]

	PIN TDB[96]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 324.015 0.25 324.115 ;
			LAYER	M2 ;
			RECT	0 324.015 0.25 324.115 ;
			LAYER	M3 ;
			RECT	0 324.015 0.25 324.115 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[96]

	PIN TDB[97]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 326.895 0.25 326.995 ;
			LAYER	M2 ;
			RECT	0 326.895 0.25 326.995 ;
			LAYER	M3 ;
			RECT	0 326.895 0.25 326.995 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[97]

	PIN TDB[98]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 329.775 0.25 329.875 ;
			LAYER	M2 ;
			RECT	0 329.775 0.25 329.875 ;
			LAYER	M3 ;
			RECT	0 329.775 0.25 329.875 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[98]

	PIN TDB[99]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 332.655 0.25 332.755 ;
			LAYER	M2 ;
			RECT	0 332.655 0.25 332.755 ;
			LAYER	M3 ;
			RECT	0 332.655 0.25 332.755 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[99]

	PIN TDB[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 27.385 0.25 27.485 ;
			LAYER	M2 ;
			RECT	0 27.385 0.25 27.485 ;
			LAYER	M3 ;
			RECT	0 27.385 0.25 27.485 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[9]

	PIN TENA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 190.45 0.25 190.55 ;
			LAYER	M2 ;
			RECT	0 190.45 0.25 190.55 ;
			LAYER	M3 ;
			RECT	0 190.45 0.25 190.55 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TENA

	PIN TENB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 224.925 0.25 225.025 ;
			LAYER	M2 ;
			RECT	0 224.925 0.25 225.025 ;
			LAYER	M3 ;
			RECT	0 224.925 0.25 225.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TENB

	PIN TWENB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 3.26 0.25 3.36 ;
			LAYER	M2 ;
			RECT	0 3.26 0.25 3.36 ;
			LAYER	M3 ;
			RECT	0 3.26 0.25 3.36 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[0]

	PIN TWENB[100]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 333.74 0.25 333.84 ;
			LAYER	M2 ;
			RECT	0 333.74 0.25 333.84 ;
			LAYER	M3 ;
			RECT	0 333.74 0.25 333.84 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[100]

	PIN TWENB[101]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 336.62 0.25 336.72 ;
			LAYER	M2 ;
			RECT	0 336.62 0.25 336.72 ;
			LAYER	M3 ;
			RECT	0 336.62 0.25 336.72 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[101]

	PIN TWENB[102]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 339.5 0.25 339.6 ;
			LAYER	M2 ;
			RECT	0 339.5 0.25 339.6 ;
			LAYER	M3 ;
			RECT	0 339.5 0.25 339.6 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[102]

	PIN TWENB[103]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 342.38 0.25 342.48 ;
			LAYER	M2 ;
			RECT	0 342.38 0.25 342.48 ;
			LAYER	M3 ;
			RECT	0 342.38 0.25 342.48 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[103]

	PIN TWENB[104]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 345.26 0.25 345.36 ;
			LAYER	M2 ;
			RECT	0 345.26 0.25 345.36 ;
			LAYER	M3 ;
			RECT	0 345.26 0.25 345.36 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[104]

	PIN TWENB[105]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 348.14 0.25 348.24 ;
			LAYER	M2 ;
			RECT	0 348.14 0.25 348.24 ;
			LAYER	M3 ;
			RECT	0 348.14 0.25 348.24 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[105]

	PIN TWENB[106]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 351.02 0.25 351.12 ;
			LAYER	M2 ;
			RECT	0 351.02 0.25 351.12 ;
			LAYER	M3 ;
			RECT	0 351.02 0.25 351.12 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[106]

	PIN TWENB[107]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 353.9 0.25 354 ;
			LAYER	M2 ;
			RECT	0 353.9 0.25 354 ;
			LAYER	M3 ;
			RECT	0 353.9 0.25 354 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[107]

	PIN TWENB[108]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 356.78 0.25 356.88 ;
			LAYER	M2 ;
			RECT	0 356.78 0.25 356.88 ;
			LAYER	M3 ;
			RECT	0 356.78 0.25 356.88 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[108]

	PIN TWENB[109]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 359.66 0.25 359.76 ;
			LAYER	M2 ;
			RECT	0 359.66 0.25 359.76 ;
			LAYER	M3 ;
			RECT	0 359.66 0.25 359.76 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[109]

	PIN TWENB[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 32.06 0.25 32.16 ;
			LAYER	M2 ;
			RECT	0 32.06 0.25 32.16 ;
			LAYER	M3 ;
			RECT	0 32.06 0.25 32.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[10]

	PIN TWENB[110]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 362.54 0.25 362.64 ;
			LAYER	M2 ;
			RECT	0 362.54 0.25 362.64 ;
			LAYER	M3 ;
			RECT	0 362.54 0.25 362.64 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[110]

	PIN TWENB[111]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 365.42 0.25 365.52 ;
			LAYER	M2 ;
			RECT	0 365.42 0.25 365.52 ;
			LAYER	M3 ;
			RECT	0 365.42 0.25 365.52 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[111]

	PIN TWENB[112]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 368.3 0.25 368.4 ;
			LAYER	M2 ;
			RECT	0 368.3 0.25 368.4 ;
			LAYER	M3 ;
			RECT	0 368.3 0.25 368.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[112]

	PIN TWENB[113]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 371.18 0.25 371.28 ;
			LAYER	M2 ;
			RECT	0 371.18 0.25 371.28 ;
			LAYER	M3 ;
			RECT	0 371.18 0.25 371.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[113]

	PIN TWENB[114]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 374.06 0.25 374.16 ;
			LAYER	M2 ;
			RECT	0 374.06 0.25 374.16 ;
			LAYER	M3 ;
			RECT	0 374.06 0.25 374.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[114]

	PIN TWENB[115]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 376.94 0.25 377.04 ;
			LAYER	M2 ;
			RECT	0 376.94 0.25 377.04 ;
			LAYER	M3 ;
			RECT	0 376.94 0.25 377.04 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[115]

	PIN TWENB[116]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 379.82 0.25 379.92 ;
			LAYER	M2 ;
			RECT	0 379.82 0.25 379.92 ;
			LAYER	M3 ;
			RECT	0 379.82 0.25 379.92 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[116]

	PIN TWENB[117]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 382.7 0.25 382.8 ;
			LAYER	M2 ;
			RECT	0 382.7 0.25 382.8 ;
			LAYER	M3 ;
			RECT	0 382.7 0.25 382.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[117]

	PIN TWENB[118]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 385.58 0.25 385.68 ;
			LAYER	M2 ;
			RECT	0 385.58 0.25 385.68 ;
			LAYER	M3 ;
			RECT	0 385.58 0.25 385.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[118]

	PIN TWENB[119]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 388.46 0.25 388.56 ;
			LAYER	M2 ;
			RECT	0 388.46 0.25 388.56 ;
			LAYER	M3 ;
			RECT	0 388.46 0.25 388.56 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[119]

	PIN TWENB[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 34.94 0.25 35.04 ;
			LAYER	M2 ;
			RECT	0 34.94 0.25 35.04 ;
			LAYER	M3 ;
			RECT	0 34.94 0.25 35.04 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[11]

	PIN TWENB[120]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 391.34 0.25 391.44 ;
			LAYER	M2 ;
			RECT	0 391.34 0.25 391.44 ;
			LAYER	M3 ;
			RECT	0 391.34 0.25 391.44 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[120]

	PIN TWENB[121]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 394.22 0.25 394.32 ;
			LAYER	M2 ;
			RECT	0 394.22 0.25 394.32 ;
			LAYER	M3 ;
			RECT	0 394.22 0.25 394.32 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[121]

	PIN TWENB[122]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 397.1 0.25 397.2 ;
			LAYER	M2 ;
			RECT	0 397.1 0.25 397.2 ;
			LAYER	M3 ;
			RECT	0 397.1 0.25 397.2 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[122]

	PIN TWENB[123]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 399.98 0.25 400.08 ;
			LAYER	M2 ;
			RECT	0 399.98 0.25 400.08 ;
			LAYER	M3 ;
			RECT	0 399.98 0.25 400.08 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[123]

	PIN TWENB[124]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 402.86 0.25 402.96 ;
			LAYER	M2 ;
			RECT	0 402.86 0.25 402.96 ;
			LAYER	M3 ;
			RECT	0 402.86 0.25 402.96 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[124]

	PIN TWENB[125]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 405.74 0.25 405.84 ;
			LAYER	M2 ;
			RECT	0 405.74 0.25 405.84 ;
			LAYER	M3 ;
			RECT	0 405.74 0.25 405.84 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[125]

	PIN TWENB[126]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 408.62 0.25 408.72 ;
			LAYER	M2 ;
			RECT	0 408.62 0.25 408.72 ;
			LAYER	M3 ;
			RECT	0 408.62 0.25 408.72 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[126]

	PIN TWENB[127]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 411.5 0.25 411.6 ;
			LAYER	M2 ;
			RECT	0 411.5 0.25 411.6 ;
			LAYER	M3 ;
			RECT	0 411.5 0.25 411.6 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[127]

	PIN TWENB[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 37.82 0.25 37.92 ;
			LAYER	M2 ;
			RECT	0 37.82 0.25 37.92 ;
			LAYER	M3 ;
			RECT	0 37.82 0.25 37.92 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[12]

	PIN TWENB[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 40.7 0.25 40.8 ;
			LAYER	M2 ;
			RECT	0 40.7 0.25 40.8 ;
			LAYER	M3 ;
			RECT	0 40.7 0.25 40.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[13]

	PIN TWENB[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 43.58 0.25 43.68 ;
			LAYER	M2 ;
			RECT	0 43.58 0.25 43.68 ;
			LAYER	M3 ;
			RECT	0 43.58 0.25 43.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[14]

	PIN TWENB[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 46.46 0.25 46.56 ;
			LAYER	M2 ;
			RECT	0 46.46 0.25 46.56 ;
			LAYER	M3 ;
			RECT	0 46.46 0.25 46.56 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[15]

	PIN TWENB[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 49.34 0.25 49.44 ;
			LAYER	M2 ;
			RECT	0 49.34 0.25 49.44 ;
			LAYER	M3 ;
			RECT	0 49.34 0.25 49.44 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[16]

	PIN TWENB[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 52.22 0.25 52.32 ;
			LAYER	M2 ;
			RECT	0 52.22 0.25 52.32 ;
			LAYER	M3 ;
			RECT	0 52.22 0.25 52.32 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[17]

	PIN TWENB[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 55.1 0.25 55.2 ;
			LAYER	M2 ;
			RECT	0 55.1 0.25 55.2 ;
			LAYER	M3 ;
			RECT	0 55.1 0.25 55.2 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[18]

	PIN TWENB[19]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 57.98 0.25 58.08 ;
			LAYER	M2 ;
			RECT	0 57.98 0.25 58.08 ;
			LAYER	M3 ;
			RECT	0 57.98 0.25 58.08 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[19]

	PIN TWENB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 6.14 0.25 6.24 ;
			LAYER	M2 ;
			RECT	0 6.14 0.25 6.24 ;
			LAYER	M3 ;
			RECT	0 6.14 0.25 6.24 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[1]

	PIN TWENB[20]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 60.86 0.25 60.96 ;
			LAYER	M2 ;
			RECT	0 60.86 0.25 60.96 ;
			LAYER	M3 ;
			RECT	0 60.86 0.25 60.96 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[20]

	PIN TWENB[21]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 63.74 0.25 63.84 ;
			LAYER	M2 ;
			RECT	0 63.74 0.25 63.84 ;
			LAYER	M3 ;
			RECT	0 63.74 0.25 63.84 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[21]

	PIN TWENB[22]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 66.62 0.25 66.72 ;
			LAYER	M2 ;
			RECT	0 66.62 0.25 66.72 ;
			LAYER	M3 ;
			RECT	0 66.62 0.25 66.72 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[22]

	PIN TWENB[23]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 69.5 0.25 69.6 ;
			LAYER	M2 ;
			RECT	0 69.5 0.25 69.6 ;
			LAYER	M3 ;
			RECT	0 69.5 0.25 69.6 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[23]

	PIN TWENB[24]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 72.38 0.25 72.48 ;
			LAYER	M2 ;
			RECT	0 72.38 0.25 72.48 ;
			LAYER	M3 ;
			RECT	0 72.38 0.25 72.48 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[24]

	PIN TWENB[25]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 75.26 0.25 75.36 ;
			LAYER	M2 ;
			RECT	0 75.26 0.25 75.36 ;
			LAYER	M3 ;
			RECT	0 75.26 0.25 75.36 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[25]

	PIN TWENB[26]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 78.14 0.25 78.24 ;
			LAYER	M2 ;
			RECT	0 78.14 0.25 78.24 ;
			LAYER	M3 ;
			RECT	0 78.14 0.25 78.24 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[26]

	PIN TWENB[27]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 81.02 0.25 81.12 ;
			LAYER	M2 ;
			RECT	0 81.02 0.25 81.12 ;
			LAYER	M3 ;
			RECT	0 81.02 0.25 81.12 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[27]

	PIN TWENB[28]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 83.9 0.25 84 ;
			LAYER	M2 ;
			RECT	0 83.9 0.25 84 ;
			LAYER	M3 ;
			RECT	0 83.9 0.25 84 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[28]

	PIN TWENB[29]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 86.78 0.25 86.88 ;
			LAYER	M2 ;
			RECT	0 86.78 0.25 86.88 ;
			LAYER	M3 ;
			RECT	0 86.78 0.25 86.88 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[29]

	PIN TWENB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 9.02 0.25 9.12 ;
			LAYER	M2 ;
			RECT	0 9.02 0.25 9.12 ;
			LAYER	M3 ;
			RECT	0 9.02 0.25 9.12 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[2]

	PIN TWENB[30]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 89.66 0.25 89.76 ;
			LAYER	M2 ;
			RECT	0 89.66 0.25 89.76 ;
			LAYER	M3 ;
			RECT	0 89.66 0.25 89.76 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[30]

	PIN TWENB[31]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 92.54 0.25 92.64 ;
			LAYER	M2 ;
			RECT	0 92.54 0.25 92.64 ;
			LAYER	M3 ;
			RECT	0 92.54 0.25 92.64 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[31]

	PIN TWENB[32]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 95.42 0.25 95.52 ;
			LAYER	M2 ;
			RECT	0 95.42 0.25 95.52 ;
			LAYER	M3 ;
			RECT	0 95.42 0.25 95.52 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[32]

	PIN TWENB[33]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 98.3 0.25 98.4 ;
			LAYER	M2 ;
			RECT	0 98.3 0.25 98.4 ;
			LAYER	M3 ;
			RECT	0 98.3 0.25 98.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[33]

	PIN TWENB[34]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 101.18 0.25 101.28 ;
			LAYER	M2 ;
			RECT	0 101.18 0.25 101.28 ;
			LAYER	M3 ;
			RECT	0 101.18 0.25 101.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[34]

	PIN TWENB[35]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 104.06 0.25 104.16 ;
			LAYER	M2 ;
			RECT	0 104.06 0.25 104.16 ;
			LAYER	M3 ;
			RECT	0 104.06 0.25 104.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[35]

	PIN TWENB[36]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 106.94 0.25 107.04 ;
			LAYER	M2 ;
			RECT	0 106.94 0.25 107.04 ;
			LAYER	M3 ;
			RECT	0 106.94 0.25 107.04 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[36]

	PIN TWENB[37]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 109.82 0.25 109.92 ;
			LAYER	M2 ;
			RECT	0 109.82 0.25 109.92 ;
			LAYER	M3 ;
			RECT	0 109.82 0.25 109.92 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[37]

	PIN TWENB[38]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 112.7 0.25 112.8 ;
			LAYER	M2 ;
			RECT	0 112.7 0.25 112.8 ;
			LAYER	M3 ;
			RECT	0 112.7 0.25 112.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[38]

	PIN TWENB[39]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 115.58 0.25 115.68 ;
			LAYER	M2 ;
			RECT	0 115.58 0.25 115.68 ;
			LAYER	M3 ;
			RECT	0 115.58 0.25 115.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[39]

	PIN TWENB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 11.9 0.25 12 ;
			LAYER	M2 ;
			RECT	0 11.9 0.25 12 ;
			LAYER	M3 ;
			RECT	0 11.9 0.25 12 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[3]

	PIN TWENB[40]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 118.46 0.25 118.56 ;
			LAYER	M2 ;
			RECT	0 118.46 0.25 118.56 ;
			LAYER	M3 ;
			RECT	0 118.46 0.25 118.56 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[40]

	PIN TWENB[41]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 121.34 0.25 121.44 ;
			LAYER	M2 ;
			RECT	0 121.34 0.25 121.44 ;
			LAYER	M3 ;
			RECT	0 121.34 0.25 121.44 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[41]

	PIN TWENB[42]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 124.22 0.25 124.32 ;
			LAYER	M2 ;
			RECT	0 124.22 0.25 124.32 ;
			LAYER	M3 ;
			RECT	0 124.22 0.25 124.32 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[42]

	PIN TWENB[43]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 127.1 0.25 127.2 ;
			LAYER	M2 ;
			RECT	0 127.1 0.25 127.2 ;
			LAYER	M3 ;
			RECT	0 127.1 0.25 127.2 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[43]

	PIN TWENB[44]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 129.98 0.25 130.08 ;
			LAYER	M2 ;
			RECT	0 129.98 0.25 130.08 ;
			LAYER	M3 ;
			RECT	0 129.98 0.25 130.08 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[44]

	PIN TWENB[45]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 132.86 0.25 132.96 ;
			LAYER	M2 ;
			RECT	0 132.86 0.25 132.96 ;
			LAYER	M3 ;
			RECT	0 132.86 0.25 132.96 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[45]

	PIN TWENB[46]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 135.74 0.25 135.84 ;
			LAYER	M2 ;
			RECT	0 135.74 0.25 135.84 ;
			LAYER	M3 ;
			RECT	0 135.74 0.25 135.84 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[46]

	PIN TWENB[47]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 138.62 0.25 138.72 ;
			LAYER	M2 ;
			RECT	0 138.62 0.25 138.72 ;
			LAYER	M3 ;
			RECT	0 138.62 0.25 138.72 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[47]

	PIN TWENB[48]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 141.5 0.25 141.6 ;
			LAYER	M2 ;
			RECT	0 141.5 0.25 141.6 ;
			LAYER	M3 ;
			RECT	0 141.5 0.25 141.6 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[48]

	PIN TWENB[49]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 144.38 0.25 144.48 ;
			LAYER	M2 ;
			RECT	0 144.38 0.25 144.48 ;
			LAYER	M3 ;
			RECT	0 144.38 0.25 144.48 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[49]

	PIN TWENB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 14.78 0.25 14.88 ;
			LAYER	M2 ;
			RECT	0 14.78 0.25 14.88 ;
			LAYER	M3 ;
			RECT	0 14.78 0.25 14.88 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[4]

	PIN TWENB[50]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 147.26 0.25 147.36 ;
			LAYER	M2 ;
			RECT	0 147.26 0.25 147.36 ;
			LAYER	M3 ;
			RECT	0 147.26 0.25 147.36 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[50]

	PIN TWENB[51]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 150.14 0.25 150.24 ;
			LAYER	M2 ;
			RECT	0 150.14 0.25 150.24 ;
			LAYER	M3 ;
			RECT	0 150.14 0.25 150.24 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[51]

	PIN TWENB[52]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 153.02 0.25 153.12 ;
			LAYER	M2 ;
			RECT	0 153.02 0.25 153.12 ;
			LAYER	M3 ;
			RECT	0 153.02 0.25 153.12 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[52]

	PIN TWENB[53]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 155.9 0.25 156 ;
			LAYER	M2 ;
			RECT	0 155.9 0.25 156 ;
			LAYER	M3 ;
			RECT	0 155.9 0.25 156 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[53]

	PIN TWENB[54]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 158.78 0.25 158.88 ;
			LAYER	M2 ;
			RECT	0 158.78 0.25 158.88 ;
			LAYER	M3 ;
			RECT	0 158.78 0.25 158.88 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[54]

	PIN TWENB[55]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 161.66 0.25 161.76 ;
			LAYER	M2 ;
			RECT	0 161.66 0.25 161.76 ;
			LAYER	M3 ;
			RECT	0 161.66 0.25 161.76 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[55]

	PIN TWENB[56]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 164.54 0.25 164.64 ;
			LAYER	M2 ;
			RECT	0 164.54 0.25 164.64 ;
			LAYER	M3 ;
			RECT	0 164.54 0.25 164.64 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[56]

	PIN TWENB[57]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 167.42 0.25 167.52 ;
			LAYER	M2 ;
			RECT	0 167.42 0.25 167.52 ;
			LAYER	M3 ;
			RECT	0 167.42 0.25 167.52 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[57]

	PIN TWENB[58]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 170.3 0.25 170.4 ;
			LAYER	M2 ;
			RECT	0 170.3 0.25 170.4 ;
			LAYER	M3 ;
			RECT	0 170.3 0.25 170.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[58]

	PIN TWENB[59]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 173.18 0.25 173.28 ;
			LAYER	M2 ;
			RECT	0 173.18 0.25 173.28 ;
			LAYER	M3 ;
			RECT	0 173.18 0.25 173.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[59]

	PIN TWENB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 17.66 0.25 17.76 ;
			LAYER	M2 ;
			RECT	0 17.66 0.25 17.76 ;
			LAYER	M3 ;
			RECT	0 17.66 0.25 17.76 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[5]

	PIN TWENB[60]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 176.06 0.25 176.16 ;
			LAYER	M2 ;
			RECT	0 176.06 0.25 176.16 ;
			LAYER	M3 ;
			RECT	0 176.06 0.25 176.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[60]

	PIN TWENB[61]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 178.94 0.25 179.04 ;
			LAYER	M2 ;
			RECT	0 178.94 0.25 179.04 ;
			LAYER	M3 ;
			RECT	0 178.94 0.25 179.04 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[61]

	PIN TWENB[62]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 181.82 0.25 181.92 ;
			LAYER	M2 ;
			RECT	0 181.82 0.25 181.92 ;
			LAYER	M3 ;
			RECT	0 181.82 0.25 181.92 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[62]

	PIN TWENB[63]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 184.7 0.25 184.8 ;
			LAYER	M2 ;
			RECT	0 184.7 0.25 184.8 ;
			LAYER	M3 ;
			RECT	0 184.7 0.25 184.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[63]

	PIN TWENB[64]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 230.06 0.25 230.16 ;
			LAYER	M2 ;
			RECT	0 230.06 0.25 230.16 ;
			LAYER	M3 ;
			RECT	0 230.06 0.25 230.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[64]

	PIN TWENB[65]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 232.94 0.25 233.04 ;
			LAYER	M2 ;
			RECT	0 232.94 0.25 233.04 ;
			LAYER	M3 ;
			RECT	0 232.94 0.25 233.04 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[65]

	PIN TWENB[66]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 235.82 0.25 235.92 ;
			LAYER	M2 ;
			RECT	0 235.82 0.25 235.92 ;
			LAYER	M3 ;
			RECT	0 235.82 0.25 235.92 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[66]

	PIN TWENB[67]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 238.7 0.25 238.8 ;
			LAYER	M2 ;
			RECT	0 238.7 0.25 238.8 ;
			LAYER	M3 ;
			RECT	0 238.7 0.25 238.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[67]

	PIN TWENB[68]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 241.58 0.25 241.68 ;
			LAYER	M2 ;
			RECT	0 241.58 0.25 241.68 ;
			LAYER	M3 ;
			RECT	0 241.58 0.25 241.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[68]

	PIN TWENB[69]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 244.46 0.25 244.56 ;
			LAYER	M2 ;
			RECT	0 244.46 0.25 244.56 ;
			LAYER	M3 ;
			RECT	0 244.46 0.25 244.56 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[69]

	PIN TWENB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 20.54 0.25 20.64 ;
			LAYER	M2 ;
			RECT	0 20.54 0.25 20.64 ;
			LAYER	M3 ;
			RECT	0 20.54 0.25 20.64 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[6]

	PIN TWENB[70]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 247.34 0.25 247.44 ;
			LAYER	M2 ;
			RECT	0 247.34 0.25 247.44 ;
			LAYER	M3 ;
			RECT	0 247.34 0.25 247.44 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[70]

	PIN TWENB[71]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 250.22 0.25 250.32 ;
			LAYER	M2 ;
			RECT	0 250.22 0.25 250.32 ;
			LAYER	M3 ;
			RECT	0 250.22 0.25 250.32 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[71]

	PIN TWENB[72]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 253.1 0.25 253.2 ;
			LAYER	M2 ;
			RECT	0 253.1 0.25 253.2 ;
			LAYER	M3 ;
			RECT	0 253.1 0.25 253.2 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[72]

	PIN TWENB[73]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 255.98 0.25 256.08 ;
			LAYER	M2 ;
			RECT	0 255.98 0.25 256.08 ;
			LAYER	M3 ;
			RECT	0 255.98 0.25 256.08 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[73]

	PIN TWENB[74]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 258.86 0.25 258.96 ;
			LAYER	M2 ;
			RECT	0 258.86 0.25 258.96 ;
			LAYER	M3 ;
			RECT	0 258.86 0.25 258.96 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[74]

	PIN TWENB[75]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 261.74 0.25 261.84 ;
			LAYER	M2 ;
			RECT	0 261.74 0.25 261.84 ;
			LAYER	M3 ;
			RECT	0 261.74 0.25 261.84 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[75]

	PIN TWENB[76]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 264.62 0.25 264.72 ;
			LAYER	M2 ;
			RECT	0 264.62 0.25 264.72 ;
			LAYER	M3 ;
			RECT	0 264.62 0.25 264.72 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[76]

	PIN TWENB[77]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 267.5 0.25 267.6 ;
			LAYER	M2 ;
			RECT	0 267.5 0.25 267.6 ;
			LAYER	M3 ;
			RECT	0 267.5 0.25 267.6 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[77]

	PIN TWENB[78]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 270.38 0.25 270.48 ;
			LAYER	M2 ;
			RECT	0 270.38 0.25 270.48 ;
			LAYER	M3 ;
			RECT	0 270.38 0.25 270.48 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[78]

	PIN TWENB[79]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 273.26 0.25 273.36 ;
			LAYER	M2 ;
			RECT	0 273.26 0.25 273.36 ;
			LAYER	M3 ;
			RECT	0 273.26 0.25 273.36 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[79]

	PIN TWENB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 23.42 0.25 23.52 ;
			LAYER	M2 ;
			RECT	0 23.42 0.25 23.52 ;
			LAYER	M3 ;
			RECT	0 23.42 0.25 23.52 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[7]

	PIN TWENB[80]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 276.14 0.25 276.24 ;
			LAYER	M2 ;
			RECT	0 276.14 0.25 276.24 ;
			LAYER	M3 ;
			RECT	0 276.14 0.25 276.24 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[80]

	PIN TWENB[81]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 279.02 0.25 279.12 ;
			LAYER	M2 ;
			RECT	0 279.02 0.25 279.12 ;
			LAYER	M3 ;
			RECT	0 279.02 0.25 279.12 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[81]

	PIN TWENB[82]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 281.9 0.25 282 ;
			LAYER	M2 ;
			RECT	0 281.9 0.25 282 ;
			LAYER	M3 ;
			RECT	0 281.9 0.25 282 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[82]

	PIN TWENB[83]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 284.78 0.25 284.88 ;
			LAYER	M2 ;
			RECT	0 284.78 0.25 284.88 ;
			LAYER	M3 ;
			RECT	0 284.78 0.25 284.88 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[83]

	PIN TWENB[84]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 287.66 0.25 287.76 ;
			LAYER	M2 ;
			RECT	0 287.66 0.25 287.76 ;
			LAYER	M3 ;
			RECT	0 287.66 0.25 287.76 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[84]

	PIN TWENB[85]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 290.54 0.25 290.64 ;
			LAYER	M2 ;
			RECT	0 290.54 0.25 290.64 ;
			LAYER	M3 ;
			RECT	0 290.54 0.25 290.64 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[85]

	PIN TWENB[86]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 293.42 0.25 293.52 ;
			LAYER	M2 ;
			RECT	0 293.42 0.25 293.52 ;
			LAYER	M3 ;
			RECT	0 293.42 0.25 293.52 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[86]

	PIN TWENB[87]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 296.3 0.25 296.4 ;
			LAYER	M2 ;
			RECT	0 296.3 0.25 296.4 ;
			LAYER	M3 ;
			RECT	0 296.3 0.25 296.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[87]

	PIN TWENB[88]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 299.18 0.25 299.28 ;
			LAYER	M2 ;
			RECT	0 299.18 0.25 299.28 ;
			LAYER	M3 ;
			RECT	0 299.18 0.25 299.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[88]

	PIN TWENB[89]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 302.06 0.25 302.16 ;
			LAYER	M2 ;
			RECT	0 302.06 0.25 302.16 ;
			LAYER	M3 ;
			RECT	0 302.06 0.25 302.16 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[89]

	PIN TWENB[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 26.3 0.25 26.4 ;
			LAYER	M2 ;
			RECT	0 26.3 0.25 26.4 ;
			LAYER	M3 ;
			RECT	0 26.3 0.25 26.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[8]

	PIN TWENB[90]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 304.94 0.25 305.04 ;
			LAYER	M2 ;
			RECT	0 304.94 0.25 305.04 ;
			LAYER	M3 ;
			RECT	0 304.94 0.25 305.04 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[90]

	PIN TWENB[91]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 307.82 0.25 307.92 ;
			LAYER	M2 ;
			RECT	0 307.82 0.25 307.92 ;
			LAYER	M3 ;
			RECT	0 307.82 0.25 307.92 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[91]

	PIN TWENB[92]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 310.7 0.25 310.8 ;
			LAYER	M2 ;
			RECT	0 310.7 0.25 310.8 ;
			LAYER	M3 ;
			RECT	0 310.7 0.25 310.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[92]

	PIN TWENB[93]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 313.58 0.25 313.68 ;
			LAYER	M2 ;
			RECT	0 313.58 0.25 313.68 ;
			LAYER	M3 ;
			RECT	0 313.58 0.25 313.68 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[93]

	PIN TWENB[94]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 316.46 0.25 316.56 ;
			LAYER	M2 ;
			RECT	0 316.46 0.25 316.56 ;
			LAYER	M3 ;
			RECT	0 316.46 0.25 316.56 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[94]

	PIN TWENB[95]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 319.34 0.25 319.44 ;
			LAYER	M2 ;
			RECT	0 319.34 0.25 319.44 ;
			LAYER	M3 ;
			RECT	0 319.34 0.25 319.44 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[95]

	PIN TWENB[96]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 322.22 0.25 322.32 ;
			LAYER	M2 ;
			RECT	0 322.22 0.25 322.32 ;
			LAYER	M3 ;
			RECT	0 322.22 0.25 322.32 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[96]

	PIN TWENB[97]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 325.1 0.25 325.2 ;
			LAYER	M2 ;
			RECT	0 325.1 0.25 325.2 ;
			LAYER	M3 ;
			RECT	0 325.1 0.25 325.2 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[97]

	PIN TWENB[98]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 327.98 0.25 328.08 ;
			LAYER	M2 ;
			RECT	0 327.98 0.25 328.08 ;
			LAYER	M3 ;
			RECT	0 327.98 0.25 328.08 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[98]

	PIN TWENB[99]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 330.86 0.25 330.96 ;
			LAYER	M2 ;
			RECT	0 330.86 0.25 330.96 ;
			LAYER	M3 ;
			RECT	0 330.86 0.25 330.96 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[99]

	PIN TWENB[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 29.18 0.25 29.28 ;
			LAYER	M2 ;
			RECT	0 29.18 0.25 29.28 ;
			LAYER	M3 ;
			RECT	0 29.18 0.25 29.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TWENB[9]

	PIN VDDCE
		USE POWER ;
		DIRECTION INOUT ;
		PORT
			LAYER	M4 ;
			RECT	0 411.415 21.975 411.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 356.695 21.975 356.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 353.815 21.975 353.965 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 408.535 21.975 408.685 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 350.935 21.975 351.085 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 348.055 21.975 348.205 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 345.175 21.975 345.325 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 342.295 21.975 342.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 339.415 21.975 339.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 336.535 21.975 336.685 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 333.655 21.975 333.805 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 330.775 21.975 330.925 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 327.895 21.975 328.045 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 325.015 21.975 325.165 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 405.655 21.975 405.805 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 322.135 21.975 322.285 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 319.255 21.975 319.405 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 316.375 21.975 316.525 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 313.495 21.975 313.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 310.615 21.975 310.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 307.735 21.975 307.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 304.855 21.975 305.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 301.975 21.975 302.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 299.095 21.975 299.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 296.215 21.975 296.365 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 402.775 21.975 402.925 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 293.335 21.975 293.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 290.455 21.975 290.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 287.575 21.975 287.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 284.695 21.975 284.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 281.815 21.975 281.965 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 278.935 21.975 279.085 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 276.055 21.975 276.205 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 273.175 21.975 273.325 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 270.295 21.975 270.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 267.415 21.975 267.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 399.895 21.975 400.045 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 264.535 21.975 264.685 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 261.655 21.975 261.805 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 258.775 21.975 258.925 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 255.895 21.975 256.045 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 253.015 21.975 253.165 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 250.135 21.975 250.285 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 247.255 21.975 247.405 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 244.375 21.975 244.525 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 241.495 21.975 241.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 238.615 21.975 238.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 397.015 21.975 397.165 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 235.735 21.975 235.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 232.855 21.975 233.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 229.975 21.975 230.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 394.135 21.975 394.285 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 184.735 21.975 184.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 181.855 21.975 182.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 178.975 21.975 179.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 176.095 21.975 176.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 391.255 21.975 391.405 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 173.215 21.975 173.365 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 170.335 21.975 170.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 167.455 21.975 167.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 164.575 21.975 164.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 161.695 21.975 161.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 158.815 21.975 158.965 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 155.935 21.975 156.085 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 153.055 21.975 153.205 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 150.175 21.975 150.325 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 147.295 21.975 147.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 388.375 21.975 388.525 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 144.415 21.975 144.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 141.535 21.975 141.685 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 138.655 21.975 138.805 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 135.775 21.975 135.925 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 132.895 21.975 133.045 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 130.015 21.975 130.165 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 127.135 21.975 127.285 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 124.255 21.975 124.405 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 121.375 21.975 121.525 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 118.495 21.975 118.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 385.495 21.975 385.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 115.615 21.975 115.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 112.735 21.975 112.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 109.855 21.975 110.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 106.975 21.975 107.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 104.095 21.975 104.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 101.215 21.975 101.365 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 98.335 21.975 98.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 95.455 21.975 95.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 92.575 21.975 92.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 89.695 21.975 89.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 382.615 21.975 382.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 86.815 21.975 86.965 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 83.935 21.975 84.085 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 81.055 21.975 81.205 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 78.175 21.975 78.325 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 75.295 21.975 75.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 72.415 21.975 72.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 69.535 21.975 69.685 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 66.655 21.975 66.805 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 63.775 21.975 63.925 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 60.895 21.975 61.045 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 379.735 21.975 379.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 58.015 21.975 58.165 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 55.135 21.975 55.285 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 52.255 21.975 52.405 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 49.375 21.975 49.525 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 46.495 21.975 46.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 43.615 21.975 43.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 40.735 21.975 40.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 37.855 21.975 38.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 34.975 21.975 35.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.095 21.975 32.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 376.855 21.975 377.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 29.215 21.975 29.365 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 26.335 21.975 26.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 23.455 21.975 23.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 20.575 21.975 20.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 17.695 21.975 17.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 14.815 21.975 14.965 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 11.935 21.975 12.085 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.055 21.975 9.205 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.175 21.975 6.325 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.295 21.975 3.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 373.975 21.975 374.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 371.095 21.975 371.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 368.215 21.975 368.365 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 365.335 21.975 365.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 362.455 21.975 362.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 359.575 21.975 359.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 191.38 21.975 191.57 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 192.36 21.975 192.55 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 195.315 21.975 195.505 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 199.25 21.975 199.44 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 200.235 21.975 200.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 203.185 21.975 203.375 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 207.12 21.975 207.31 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 207.615 21.975 207.805 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 211.55 21.975 211.74 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 214.505 21.975 214.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 215.485 21.975 215.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 219.425 21.975 219.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 222.375 21.975 222.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 223.325 21.975 223.515 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 187.095 21.975 187.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 227.615 21.975 227.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 414.295 21.975 414.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.415 21.975 0.565 ;
		END

	END VDDCE

	PIN VDDPE
		USE POWER ;
		DIRECTION INOUT ;
		PORT
			LAYER	M4 ;
			RECT	0 188.425 21.975 188.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 190.43 21.975 190.62 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 193.345 21.975 193.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 194.33 21.975 194.52 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 196.3 21.975 196.49 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 197.28 21.975 197.47 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 198.265 21.975 198.455 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 201.22 21.975 201.41 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 205.155 21.975 205.345 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 206.14 21.975 206.33 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 208.6 21.975 208.79 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 209.58 21.975 209.77 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 213.52 21.975 213.71 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 216.47 21.975 216.66 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 217.455 21.975 217.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 218.44 21.975 218.63 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 220.405 21.975 220.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 221.39 21.975 221.58 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 224.31 21.975 224.5 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 226.31 21.975 226.5 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 413.835 21.975 413.985 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 356.235 21.975 356.385 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 353.355 21.975 353.505 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 350.475 21.975 350.625 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 347.595 21.975 347.745 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 344.715 21.975 344.865 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 341.835 21.975 341.985 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 408.075 21.975 408.225 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 338.955 21.975 339.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 336.075 21.975 336.225 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 333.195 21.975 333.345 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 330.315 21.975 330.465 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 327.435 21.975 327.585 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 324.555 21.975 324.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 321.675 21.975 321.825 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 318.795 21.975 318.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 315.915 21.975 316.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 313.035 21.975 313.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 405.195 21.975 405.345 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 310.155 21.975 310.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 307.275 21.975 307.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 304.395 21.975 304.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 301.515 21.975 301.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 298.635 21.975 298.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 295.755 21.975 295.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 292.875 21.975 293.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 289.995 21.975 290.145 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 287.115 21.975 287.265 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 284.235 21.975 284.385 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 402.315 21.975 402.465 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 281.355 21.975 281.505 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 278.475 21.975 278.625 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 275.595 21.975 275.745 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 272.715 21.975 272.865 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 269.835 21.975 269.985 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 266.955 21.975 267.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 264.075 21.975 264.225 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 261.195 21.975 261.345 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 258.315 21.975 258.465 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 255.435 21.975 255.585 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 399.435 21.975 399.585 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 252.555 21.975 252.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 249.675 21.975 249.825 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 246.795 21.975 246.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 243.915 21.975 244.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 241.035 21.975 241.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 238.155 21.975 238.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 235.275 21.975 235.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 232.395 21.975 232.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 396.555 21.975 396.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 393.675 21.975 393.825 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 182.315 21.975 182.465 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 179.435 21.975 179.585 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 176.555 21.975 176.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 173.675 21.975 173.825 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 170.795 21.975 170.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 167.915 21.975 168.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 165.035 21.975 165.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 162.155 21.975 162.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 390.795 21.975 390.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 159.275 21.975 159.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 156.395 21.975 156.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 153.515 21.975 153.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 150.635 21.975 150.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 147.755 21.975 147.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 144.875 21.975 145.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 141.995 21.975 142.145 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 139.115 21.975 139.265 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 136.235 21.975 136.385 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 133.355 21.975 133.505 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 387.915 21.975 388.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 130.475 21.975 130.625 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 127.595 21.975 127.745 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 124.715 21.975 124.865 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 121.835 21.975 121.985 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 118.955 21.975 119.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 116.075 21.975 116.225 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 113.195 21.975 113.345 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 110.315 21.975 110.465 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 107.435 21.975 107.585 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 104.555 21.975 104.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 385.035 21.975 385.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 101.675 21.975 101.825 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 98.795 21.975 98.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 95.915 21.975 96.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 93.035 21.975 93.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 90.155 21.975 90.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 87.275 21.975 87.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 84.395 21.975 84.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 81.515 21.975 81.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 78.635 21.975 78.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 75.755 21.975 75.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 382.155 21.975 382.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 72.875 21.975 73.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 69.995 21.975 70.145 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 67.115 21.975 67.265 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 64.235 21.975 64.385 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 61.355 21.975 61.505 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 58.475 21.975 58.625 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 55.595 21.975 55.745 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 52.715 21.975 52.865 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 49.835 21.975 49.985 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 46.955 21.975 47.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 379.275 21.975 379.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 44.075 21.975 44.225 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 41.195 21.975 41.345 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 38.315 21.975 38.465 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 35.435 21.975 35.585 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.555 21.975 32.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 29.675 21.975 29.825 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 26.795 21.975 26.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 23.915 21.975 24.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 21.035 21.975 21.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 18.155 21.975 18.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 376.395 21.975 376.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 15.275 21.975 15.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 12.395 21.975 12.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.515 21.975 9.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.635 21.975 6.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.755 21.975 3.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.875 21.975 1.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 373.515 21.975 373.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 370.635 21.975 370.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 410.955 21.975 411.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 367.755 21.975 367.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 364.875 21.975 365.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 361.995 21.975 362.145 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 359.115 21.975 359.265 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 414.525 21.975 414.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.185 21.975 0.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 186.635 21.975 186.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 228.075 21.975 228.225 ;
		END

	END VDDPE

	PIN VSSE
		USE GROUND ;
		DIRECTION INOUT ;
		PORT
			LAYER	M4 ;
			RECT	0 414.065 21.975 414.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.645 21.975 0.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 186.865 21.975 187.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 227.845 21.975 227.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 411.185 21.975 411.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 356.465 21.975 356.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 353.585 21.975 353.735 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 350.705 21.975 350.855 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 347.825 21.975 347.975 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 408.305 21.975 408.455 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 344.945 21.975 345.095 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 342.065 21.975 342.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 339.185 21.975 339.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 336.305 21.975 336.455 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 333.425 21.975 333.575 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 330.545 21.975 330.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 327.665 21.975 327.815 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 324.785 21.975 324.935 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 321.905 21.975 322.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 319.025 21.975 319.175 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 405.425 21.975 405.575 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 316.145 21.975 316.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 313.265 21.975 313.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 310.385 21.975 310.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 307.505 21.975 307.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 304.625 21.975 304.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 301.745 21.975 301.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 298.865 21.975 299.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 295.985 21.975 296.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 293.105 21.975 293.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 290.225 21.975 290.375 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 402.545 21.975 402.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 287.345 21.975 287.495 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 284.465 21.975 284.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 281.585 21.975 281.735 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 278.705 21.975 278.855 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 275.825 21.975 275.975 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 272.945 21.975 273.095 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 270.065 21.975 270.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 267.185 21.975 267.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 264.305 21.975 264.455 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 261.425 21.975 261.575 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 399.665 21.975 399.815 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 258.545 21.975 258.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 255.665 21.975 255.815 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 252.785 21.975 252.935 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 249.905 21.975 250.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 247.025 21.975 247.175 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 244.145 21.975 244.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 241.265 21.975 241.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 238.385 21.975 238.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 235.505 21.975 235.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 232.625 21.975 232.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 396.785 21.975 396.935 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 229.745 21.975 229.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 393.905 21.975 394.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 184.965 21.975 185.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 182.085 21.975 182.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 179.205 21.975 179.355 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 176.325 21.975 176.475 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 173.445 21.975 173.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 170.565 21.975 170.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 167.685 21.975 167.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 391.025 21.975 391.175 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 164.805 21.975 164.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 161.925 21.975 162.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 159.045 21.975 159.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 156.165 21.975 156.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 153.285 21.975 153.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 150.405 21.975 150.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 147.525 21.975 147.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 144.645 21.975 144.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 141.765 21.975 141.915 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 138.885 21.975 139.035 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 388.145 21.975 388.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 136.005 21.975 136.155 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 133.125 21.975 133.275 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 130.245 21.975 130.395 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 127.365 21.975 127.515 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 124.485 21.975 124.635 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 121.605 21.975 121.755 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 118.725 21.975 118.875 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 115.845 21.975 115.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 112.965 21.975 113.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 110.085 21.975 110.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 385.265 21.975 385.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 107.205 21.975 107.355 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 104.325 21.975 104.475 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 101.445 21.975 101.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 98.565 21.975 98.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 95.685 21.975 95.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 92.805 21.975 92.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 89.925 21.975 90.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 87.045 21.975 87.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 84.165 21.975 84.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 81.285 21.975 81.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 382.385 21.975 382.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 78.405 21.975 78.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 75.525 21.975 75.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 72.645 21.975 72.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 69.765 21.975 69.915 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 66.885 21.975 67.035 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 64.005 21.975 64.155 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 61.125 21.975 61.275 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 58.245 21.975 58.395 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 55.365 21.975 55.515 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 52.485 21.975 52.635 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 379.505 21.975 379.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 49.605 21.975 49.755 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 46.725 21.975 46.875 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 43.845 21.975 43.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 40.965 21.975 41.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 38.085 21.975 38.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 35.205 21.975 35.355 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.325 21.975 32.475 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 29.445 21.975 29.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 26.565 21.975 26.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 23.685 21.975 23.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 376.625 21.975 376.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 20.805 21.975 20.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 17.925 21.975 18.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 15.045 21.975 15.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 12.165 21.975 12.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.285 21.975 9.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.405 21.975 6.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.525 21.975 3.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 373.745 21.975 373.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 370.865 21.975 371.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 367.985 21.975 368.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 365.105 21.975 365.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 362.225 21.975 362.375 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 359.345 21.975 359.495 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 413.605 21.975 413.755 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 187.935 21.975 188.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 188.915 21.975 189.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 190.885 21.975 191.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 356.005 21.975 356.155 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 353.125 21.975 353.275 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 350.245 21.975 350.395 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 347.365 21.975 347.515 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 344.485 21.975 344.635 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 341.605 21.975 341.755 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 338.725 21.975 338.875 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 335.845 21.975 335.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 407.845 21.975 407.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 332.965 21.975 333.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 330.085 21.975 330.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 327.205 21.975 327.355 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 324.325 21.975 324.475 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 321.445 21.975 321.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 318.565 21.975 318.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 315.685 21.975 315.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 312.805 21.975 312.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 309.925 21.975 310.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 307.045 21.975 307.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 404.965 21.975 405.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 304.165 21.975 304.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 301.285 21.975 301.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 298.405 21.975 298.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 295.525 21.975 295.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 292.645 21.975 292.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 289.765 21.975 289.915 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 286.885 21.975 287.035 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 284.005 21.975 284.155 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 281.125 21.975 281.275 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 278.245 21.975 278.395 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 402.085 21.975 402.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 275.365 21.975 275.515 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 272.485 21.975 272.635 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 269.605 21.975 269.755 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 266.725 21.975 266.875 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 263.845 21.975 263.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 260.965 21.975 261.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 258.085 21.975 258.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 255.205 21.975 255.355 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 252.325 21.975 252.475 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 249.445 21.975 249.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 399.205 21.975 399.355 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 246.565 21.975 246.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 243.685 21.975 243.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 240.805 21.975 240.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 237.925 21.975 238.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 235.045 21.975 235.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 232.165 21.975 232.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 396.325 21.975 396.475 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 393.445 21.975 393.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 182.545 21.975 182.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 179.665 21.975 179.815 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 176.785 21.975 176.935 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 173.905 21.975 174.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 171.025 21.975 171.175 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 168.145 21.975 168.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 165.265 21.975 165.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 162.385 21.975 162.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 159.505 21.975 159.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 156.625 21.975 156.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 390.565 21.975 390.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 153.745 21.975 153.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 150.865 21.975 151.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 147.985 21.975 148.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 145.105 21.975 145.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 142.225 21.975 142.375 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 139.345 21.975 139.495 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 136.465 21.975 136.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 133.585 21.975 133.735 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 130.705 21.975 130.855 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 127.825 21.975 127.975 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 387.685 21.975 387.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 124.945 21.975 125.095 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 122.065 21.975 122.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 119.185 21.975 119.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 116.305 21.975 116.455 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 113.425 21.975 113.575 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 110.545 21.975 110.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 107.665 21.975 107.815 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 104.785 21.975 104.935 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 101.905 21.975 102.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 99.025 21.975 99.175 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 384.805 21.975 384.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 96.145 21.975 96.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 93.265 21.975 93.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 90.385 21.975 90.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 87.505 21.975 87.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 84.625 21.975 84.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 81.745 21.975 81.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 78.865 21.975 79.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 75.985 21.975 76.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 73.105 21.975 73.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 70.225 21.975 70.375 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 381.925 21.975 382.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 67.345 21.975 67.495 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 64.465 21.975 64.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 61.585 21.975 61.735 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 58.705 21.975 58.855 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 55.825 21.975 55.975 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 52.945 21.975 53.095 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 50.065 21.975 50.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 47.185 21.975 47.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 44.305 21.975 44.455 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 41.425 21.975 41.575 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 379.045 21.975 379.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 38.545 21.975 38.695 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 35.665 21.975 35.815 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.785 21.975 32.935 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 29.905 21.975 30.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 27.025 21.975 27.175 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 24.145 21.975 24.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 21.265 21.975 21.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 18.385 21.975 18.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 15.505 21.975 15.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 12.625 21.975 12.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 376.165 21.975 376.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.745 21.975 9.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.865 21.975 7.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.985 21.975 4.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 1.105 21.975 1.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 373.285 21.975 373.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 370.405 21.975 370.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 367.525 21.975 367.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 364.645 21.975 364.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 410.725 21.975 410.875 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 361.765 21.975 361.915 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 358.885 21.975 359.035 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 191.87 21.975 192.06 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 194.825 21.975 195.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 195.805 21.975 195.995 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 196.79 21.975 196.98 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 198.76 21.975 198.95 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 199.73 21.975 199.94 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 200.725 21.975 200.915 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 202.7 21.975 202.89 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 203.68 21.975 203.87 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 206.63 21.975 206.82 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 208.105 21.975 208.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 211.055 21.975 211.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 212.045 21.975 212.235 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 214.01 21.975 214.2 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 214.985 21.975 215.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 215.98 21.975 216.17 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 217.945 21.975 218.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 218.93 21.975 219.12 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 219.915 21.975 220.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 222.855 21.975 223.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 223.85 21.975 224.04 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 225.82 21.975 226.01 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 226.805 21.975 226.995 ;
		END

	END VSSE

	PIN WENB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 1.995 0.25 2.095 ;
			LAYER	M2 ;
			RECT	0 1.995 0.25 2.095 ;
			LAYER	M3 ;
			RECT	0 1.995 0.25 2.095 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[0]

	PIN WENB[100]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 335.005 0.25 335.105 ;
			LAYER	M2 ;
			RECT	0 335.005 0.25 335.105 ;
			LAYER	M3 ;
			RECT	0 335.005 0.25 335.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[100]

	PIN WENB[101]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 337.885 0.25 337.985 ;
			LAYER	M2 ;
			RECT	0 337.885 0.25 337.985 ;
			LAYER	M3 ;
			RECT	0 337.885 0.25 337.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[101]

	PIN WENB[102]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 340.765 0.25 340.865 ;
			LAYER	M2 ;
			RECT	0 340.765 0.25 340.865 ;
			LAYER	M3 ;
			RECT	0 340.765 0.25 340.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[102]

	PIN WENB[103]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 343.645 0.25 343.745 ;
			LAYER	M2 ;
			RECT	0 343.645 0.25 343.745 ;
			LAYER	M3 ;
			RECT	0 343.645 0.25 343.745 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[103]

	PIN WENB[104]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 346.525 0.25 346.625 ;
			LAYER	M2 ;
			RECT	0 346.525 0.25 346.625 ;
			LAYER	M3 ;
			RECT	0 346.525 0.25 346.625 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[104]

	PIN WENB[105]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 349.405 0.25 349.505 ;
			LAYER	M2 ;
			RECT	0 349.405 0.25 349.505 ;
			LAYER	M3 ;
			RECT	0 349.405 0.25 349.505 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[105]

	PIN WENB[106]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 352.285 0.25 352.385 ;
			LAYER	M2 ;
			RECT	0 352.285 0.25 352.385 ;
			LAYER	M3 ;
			RECT	0 352.285 0.25 352.385 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[106]

	PIN WENB[107]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 355.165 0.25 355.265 ;
			LAYER	M2 ;
			RECT	0 355.165 0.25 355.265 ;
			LAYER	M3 ;
			RECT	0 355.165 0.25 355.265 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[107]

	PIN WENB[108]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 358.045 0.25 358.145 ;
			LAYER	M2 ;
			RECT	0 358.045 0.25 358.145 ;
			LAYER	M3 ;
			RECT	0 358.045 0.25 358.145 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[108]

	PIN WENB[109]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 360.925 0.25 361.025 ;
			LAYER	M2 ;
			RECT	0 360.925 0.25 361.025 ;
			LAYER	M3 ;
			RECT	0 360.925 0.25 361.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[109]

	PIN WENB[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 30.795 0.25 30.895 ;
			LAYER	M2 ;
			RECT	0 30.795 0.25 30.895 ;
			LAYER	M3 ;
			RECT	0 30.795 0.25 30.895 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[10]

	PIN WENB[110]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 363.805 0.25 363.905 ;
			LAYER	M2 ;
			RECT	0 363.805 0.25 363.905 ;
			LAYER	M3 ;
			RECT	0 363.805 0.25 363.905 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[110]

	PIN WENB[111]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 366.685 0.25 366.785 ;
			LAYER	M2 ;
			RECT	0 366.685 0.25 366.785 ;
			LAYER	M3 ;
			RECT	0 366.685 0.25 366.785 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[111]

	PIN WENB[112]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 369.565 0.25 369.665 ;
			LAYER	M2 ;
			RECT	0 369.565 0.25 369.665 ;
			LAYER	M3 ;
			RECT	0 369.565 0.25 369.665 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[112]

	PIN WENB[113]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 372.445 0.25 372.545 ;
			LAYER	M2 ;
			RECT	0 372.445 0.25 372.545 ;
			LAYER	M3 ;
			RECT	0 372.445 0.25 372.545 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[113]

	PIN WENB[114]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 375.325 0.25 375.425 ;
			LAYER	M2 ;
			RECT	0 375.325 0.25 375.425 ;
			LAYER	M3 ;
			RECT	0 375.325 0.25 375.425 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[114]

	PIN WENB[115]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 378.205 0.25 378.305 ;
			LAYER	M2 ;
			RECT	0 378.205 0.25 378.305 ;
			LAYER	M3 ;
			RECT	0 378.205 0.25 378.305 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[115]

	PIN WENB[116]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 381.085 0.25 381.185 ;
			LAYER	M2 ;
			RECT	0 381.085 0.25 381.185 ;
			LAYER	M3 ;
			RECT	0 381.085 0.25 381.185 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[116]

	PIN WENB[117]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 383.965 0.25 384.065 ;
			LAYER	M2 ;
			RECT	0 383.965 0.25 384.065 ;
			LAYER	M3 ;
			RECT	0 383.965 0.25 384.065 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[117]

	PIN WENB[118]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 386.845 0.25 386.945 ;
			LAYER	M2 ;
			RECT	0 386.845 0.25 386.945 ;
			LAYER	M3 ;
			RECT	0 386.845 0.25 386.945 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[118]

	PIN WENB[119]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 389.725 0.25 389.825 ;
			LAYER	M2 ;
			RECT	0 389.725 0.25 389.825 ;
			LAYER	M3 ;
			RECT	0 389.725 0.25 389.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[119]

	PIN WENB[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 33.675 0.25 33.775 ;
			LAYER	M2 ;
			RECT	0 33.675 0.25 33.775 ;
			LAYER	M3 ;
			RECT	0 33.675 0.25 33.775 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[11]

	PIN WENB[120]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 392.605 0.25 392.705 ;
			LAYER	M2 ;
			RECT	0 392.605 0.25 392.705 ;
			LAYER	M3 ;
			RECT	0 392.605 0.25 392.705 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[120]

	PIN WENB[121]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 395.485 0.25 395.585 ;
			LAYER	M2 ;
			RECT	0 395.485 0.25 395.585 ;
			LAYER	M3 ;
			RECT	0 395.485 0.25 395.585 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[121]

	PIN WENB[122]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 398.365 0.25 398.465 ;
			LAYER	M2 ;
			RECT	0 398.365 0.25 398.465 ;
			LAYER	M3 ;
			RECT	0 398.365 0.25 398.465 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[122]

	PIN WENB[123]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 401.245 0.25 401.345 ;
			LAYER	M2 ;
			RECT	0 401.245 0.25 401.345 ;
			LAYER	M3 ;
			RECT	0 401.245 0.25 401.345 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[123]

	PIN WENB[124]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 404.125 0.25 404.225 ;
			LAYER	M2 ;
			RECT	0 404.125 0.25 404.225 ;
			LAYER	M3 ;
			RECT	0 404.125 0.25 404.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[124]

	PIN WENB[125]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 407.005 0.25 407.105 ;
			LAYER	M2 ;
			RECT	0 407.005 0.25 407.105 ;
			LAYER	M3 ;
			RECT	0 407.005 0.25 407.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[125]

	PIN WENB[126]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 409.885 0.25 409.985 ;
			LAYER	M2 ;
			RECT	0 409.885 0.25 409.985 ;
			LAYER	M3 ;
			RECT	0 409.885 0.25 409.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[126]

	PIN WENB[127]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 412.765 0.25 412.865 ;
			LAYER	M2 ;
			RECT	0 412.765 0.25 412.865 ;
			LAYER	M3 ;
			RECT	0 412.765 0.25 412.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[127]

	PIN WENB[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 36.555 0.25 36.655 ;
			LAYER	M2 ;
			RECT	0 36.555 0.25 36.655 ;
			LAYER	M3 ;
			RECT	0 36.555 0.25 36.655 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[12]

	PIN WENB[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 39.435 0.25 39.535 ;
			LAYER	M2 ;
			RECT	0 39.435 0.25 39.535 ;
			LAYER	M3 ;
			RECT	0 39.435 0.25 39.535 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[13]

	PIN WENB[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 42.315 0.25 42.415 ;
			LAYER	M2 ;
			RECT	0 42.315 0.25 42.415 ;
			LAYER	M3 ;
			RECT	0 42.315 0.25 42.415 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[14]

	PIN WENB[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 45.195 0.25 45.295 ;
			LAYER	M2 ;
			RECT	0 45.195 0.25 45.295 ;
			LAYER	M3 ;
			RECT	0 45.195 0.25 45.295 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[15]

	PIN WENB[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 48.075 0.25 48.175 ;
			LAYER	M2 ;
			RECT	0 48.075 0.25 48.175 ;
			LAYER	M3 ;
			RECT	0 48.075 0.25 48.175 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[16]

	PIN WENB[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 50.955 0.25 51.055 ;
			LAYER	M2 ;
			RECT	0 50.955 0.25 51.055 ;
			LAYER	M3 ;
			RECT	0 50.955 0.25 51.055 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[17]

	PIN WENB[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 53.835 0.25 53.935 ;
			LAYER	M2 ;
			RECT	0 53.835 0.25 53.935 ;
			LAYER	M3 ;
			RECT	0 53.835 0.25 53.935 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[18]

	PIN WENB[19]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 56.715 0.25 56.815 ;
			LAYER	M2 ;
			RECT	0 56.715 0.25 56.815 ;
			LAYER	M3 ;
			RECT	0 56.715 0.25 56.815 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[19]

	PIN WENB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 4.875 0.25 4.975 ;
			LAYER	M2 ;
			RECT	0 4.875 0.25 4.975 ;
			LAYER	M3 ;
			RECT	0 4.875 0.25 4.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[1]

	PIN WENB[20]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 59.595 0.25 59.695 ;
			LAYER	M2 ;
			RECT	0 59.595 0.25 59.695 ;
			LAYER	M3 ;
			RECT	0 59.595 0.25 59.695 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[20]

	PIN WENB[21]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 62.475 0.25 62.575 ;
			LAYER	M2 ;
			RECT	0 62.475 0.25 62.575 ;
			LAYER	M3 ;
			RECT	0 62.475 0.25 62.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[21]

	PIN WENB[22]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 65.355 0.25 65.455 ;
			LAYER	M2 ;
			RECT	0 65.355 0.25 65.455 ;
			LAYER	M3 ;
			RECT	0 65.355 0.25 65.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[22]

	PIN WENB[23]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 68.235 0.25 68.335 ;
			LAYER	M2 ;
			RECT	0 68.235 0.25 68.335 ;
			LAYER	M3 ;
			RECT	0 68.235 0.25 68.335 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[23]

	PIN WENB[24]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 71.115 0.25 71.215 ;
			LAYER	M2 ;
			RECT	0 71.115 0.25 71.215 ;
			LAYER	M3 ;
			RECT	0 71.115 0.25 71.215 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[24]

	PIN WENB[25]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 73.995 0.25 74.095 ;
			LAYER	M2 ;
			RECT	0 73.995 0.25 74.095 ;
			LAYER	M3 ;
			RECT	0 73.995 0.25 74.095 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[25]

	PIN WENB[26]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 76.875 0.25 76.975 ;
			LAYER	M2 ;
			RECT	0 76.875 0.25 76.975 ;
			LAYER	M3 ;
			RECT	0 76.875 0.25 76.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[26]

	PIN WENB[27]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 79.755 0.25 79.855 ;
			LAYER	M2 ;
			RECT	0 79.755 0.25 79.855 ;
			LAYER	M3 ;
			RECT	0 79.755 0.25 79.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[27]

	PIN WENB[28]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 82.635 0.25 82.735 ;
			LAYER	M2 ;
			RECT	0 82.635 0.25 82.735 ;
			LAYER	M3 ;
			RECT	0 82.635 0.25 82.735 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[28]

	PIN WENB[29]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 85.515 0.25 85.615 ;
			LAYER	M2 ;
			RECT	0 85.515 0.25 85.615 ;
			LAYER	M3 ;
			RECT	0 85.515 0.25 85.615 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[29]

	PIN WENB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 7.755 0.25 7.855 ;
			LAYER	M2 ;
			RECT	0 7.755 0.25 7.855 ;
			LAYER	M3 ;
			RECT	0 7.755 0.25 7.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[2]

	PIN WENB[30]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 88.395 0.25 88.495 ;
			LAYER	M2 ;
			RECT	0 88.395 0.25 88.495 ;
			LAYER	M3 ;
			RECT	0 88.395 0.25 88.495 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[30]

	PIN WENB[31]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 91.275 0.25 91.375 ;
			LAYER	M2 ;
			RECT	0 91.275 0.25 91.375 ;
			LAYER	M3 ;
			RECT	0 91.275 0.25 91.375 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[31]

	PIN WENB[32]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 94.155 0.25 94.255 ;
			LAYER	M2 ;
			RECT	0 94.155 0.25 94.255 ;
			LAYER	M3 ;
			RECT	0 94.155 0.25 94.255 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[32]

	PIN WENB[33]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 97.035 0.25 97.135 ;
			LAYER	M2 ;
			RECT	0 97.035 0.25 97.135 ;
			LAYER	M3 ;
			RECT	0 97.035 0.25 97.135 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[33]

	PIN WENB[34]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 99.915 0.25 100.015 ;
			LAYER	M2 ;
			RECT	0 99.915 0.25 100.015 ;
			LAYER	M3 ;
			RECT	0 99.915 0.25 100.015 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[34]

	PIN WENB[35]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 102.795 0.25 102.895 ;
			LAYER	M2 ;
			RECT	0 102.795 0.25 102.895 ;
			LAYER	M3 ;
			RECT	0 102.795 0.25 102.895 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[35]

	PIN WENB[36]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 105.675 0.25 105.775 ;
			LAYER	M2 ;
			RECT	0 105.675 0.25 105.775 ;
			LAYER	M3 ;
			RECT	0 105.675 0.25 105.775 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[36]

	PIN WENB[37]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 108.555 0.25 108.655 ;
			LAYER	M2 ;
			RECT	0 108.555 0.25 108.655 ;
			LAYER	M3 ;
			RECT	0 108.555 0.25 108.655 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[37]

	PIN WENB[38]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 111.435 0.25 111.535 ;
			LAYER	M2 ;
			RECT	0 111.435 0.25 111.535 ;
			LAYER	M3 ;
			RECT	0 111.435 0.25 111.535 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[38]

	PIN WENB[39]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 114.315 0.25 114.415 ;
			LAYER	M2 ;
			RECT	0 114.315 0.25 114.415 ;
			LAYER	M3 ;
			RECT	0 114.315 0.25 114.415 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[39]

	PIN WENB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 10.635 0.25 10.735 ;
			LAYER	M2 ;
			RECT	0 10.635 0.25 10.735 ;
			LAYER	M3 ;
			RECT	0 10.635 0.25 10.735 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[3]

	PIN WENB[40]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 117.195 0.25 117.295 ;
			LAYER	M2 ;
			RECT	0 117.195 0.25 117.295 ;
			LAYER	M3 ;
			RECT	0 117.195 0.25 117.295 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[40]

	PIN WENB[41]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 120.075 0.25 120.175 ;
			LAYER	M2 ;
			RECT	0 120.075 0.25 120.175 ;
			LAYER	M3 ;
			RECT	0 120.075 0.25 120.175 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[41]

	PIN WENB[42]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 122.955 0.25 123.055 ;
			LAYER	M2 ;
			RECT	0 122.955 0.25 123.055 ;
			LAYER	M3 ;
			RECT	0 122.955 0.25 123.055 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[42]

	PIN WENB[43]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 125.835 0.25 125.935 ;
			LAYER	M2 ;
			RECT	0 125.835 0.25 125.935 ;
			LAYER	M3 ;
			RECT	0 125.835 0.25 125.935 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[43]

	PIN WENB[44]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 128.715 0.25 128.815 ;
			LAYER	M2 ;
			RECT	0 128.715 0.25 128.815 ;
			LAYER	M3 ;
			RECT	0 128.715 0.25 128.815 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[44]

	PIN WENB[45]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 131.595 0.25 131.695 ;
			LAYER	M2 ;
			RECT	0 131.595 0.25 131.695 ;
			LAYER	M3 ;
			RECT	0 131.595 0.25 131.695 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[45]

	PIN WENB[46]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 134.475 0.25 134.575 ;
			LAYER	M2 ;
			RECT	0 134.475 0.25 134.575 ;
			LAYER	M3 ;
			RECT	0 134.475 0.25 134.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[46]

	PIN WENB[47]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 137.355 0.25 137.455 ;
			LAYER	M2 ;
			RECT	0 137.355 0.25 137.455 ;
			LAYER	M3 ;
			RECT	0 137.355 0.25 137.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[47]

	PIN WENB[48]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 140.235 0.25 140.335 ;
			LAYER	M2 ;
			RECT	0 140.235 0.25 140.335 ;
			LAYER	M3 ;
			RECT	0 140.235 0.25 140.335 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[48]

	PIN WENB[49]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 143.115 0.25 143.215 ;
			LAYER	M2 ;
			RECT	0 143.115 0.25 143.215 ;
			LAYER	M3 ;
			RECT	0 143.115 0.25 143.215 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[49]

	PIN WENB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 13.515 0.25 13.615 ;
			LAYER	M2 ;
			RECT	0 13.515 0.25 13.615 ;
			LAYER	M3 ;
			RECT	0 13.515 0.25 13.615 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[4]

	PIN WENB[50]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 145.995 0.25 146.095 ;
			LAYER	M2 ;
			RECT	0 145.995 0.25 146.095 ;
			LAYER	M3 ;
			RECT	0 145.995 0.25 146.095 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[50]

	PIN WENB[51]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 148.875 0.25 148.975 ;
			LAYER	M2 ;
			RECT	0 148.875 0.25 148.975 ;
			LAYER	M3 ;
			RECT	0 148.875 0.25 148.975 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[51]

	PIN WENB[52]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 151.755 0.25 151.855 ;
			LAYER	M2 ;
			RECT	0 151.755 0.25 151.855 ;
			LAYER	M3 ;
			RECT	0 151.755 0.25 151.855 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[52]

	PIN WENB[53]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 154.635 0.25 154.735 ;
			LAYER	M2 ;
			RECT	0 154.635 0.25 154.735 ;
			LAYER	M3 ;
			RECT	0 154.635 0.25 154.735 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[53]

	PIN WENB[54]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 157.515 0.25 157.615 ;
			LAYER	M2 ;
			RECT	0 157.515 0.25 157.615 ;
			LAYER	M3 ;
			RECT	0 157.515 0.25 157.615 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[54]

	PIN WENB[55]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 160.395 0.25 160.495 ;
			LAYER	M2 ;
			RECT	0 160.395 0.25 160.495 ;
			LAYER	M3 ;
			RECT	0 160.395 0.25 160.495 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[55]

	PIN WENB[56]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 163.275 0.25 163.375 ;
			LAYER	M2 ;
			RECT	0 163.275 0.25 163.375 ;
			LAYER	M3 ;
			RECT	0 163.275 0.25 163.375 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[56]

	PIN WENB[57]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 166.155 0.25 166.255 ;
			LAYER	M2 ;
			RECT	0 166.155 0.25 166.255 ;
			LAYER	M3 ;
			RECT	0 166.155 0.25 166.255 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[57]

	PIN WENB[58]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 169.035 0.25 169.135 ;
			LAYER	M2 ;
			RECT	0 169.035 0.25 169.135 ;
			LAYER	M3 ;
			RECT	0 169.035 0.25 169.135 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[58]

	PIN WENB[59]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 171.915 0.25 172.015 ;
			LAYER	M2 ;
			RECT	0 171.915 0.25 172.015 ;
			LAYER	M3 ;
			RECT	0 171.915 0.25 172.015 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[59]

	PIN WENB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 16.395 0.25 16.495 ;
			LAYER	M2 ;
			RECT	0 16.395 0.25 16.495 ;
			LAYER	M3 ;
			RECT	0 16.395 0.25 16.495 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[5]

	PIN WENB[60]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 174.795 0.25 174.895 ;
			LAYER	M2 ;
			RECT	0 174.795 0.25 174.895 ;
			LAYER	M3 ;
			RECT	0 174.795 0.25 174.895 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[60]

	PIN WENB[61]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 177.675 0.25 177.775 ;
			LAYER	M2 ;
			RECT	0 177.675 0.25 177.775 ;
			LAYER	M3 ;
			RECT	0 177.675 0.25 177.775 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[61]

	PIN WENB[62]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 180.555 0.25 180.655 ;
			LAYER	M2 ;
			RECT	0 180.555 0.25 180.655 ;
			LAYER	M3 ;
			RECT	0 180.555 0.25 180.655 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[62]

	PIN WENB[63]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 183.435 0.25 183.535 ;
			LAYER	M2 ;
			RECT	0 183.435 0.25 183.535 ;
			LAYER	M3 ;
			RECT	0 183.435 0.25 183.535 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[63]

	PIN WENB[64]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 231.325 0.25 231.425 ;
			LAYER	M2 ;
			RECT	0 231.325 0.25 231.425 ;
			LAYER	M3 ;
			RECT	0 231.325 0.25 231.425 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[64]

	PIN WENB[65]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 234.205 0.25 234.305 ;
			LAYER	M2 ;
			RECT	0 234.205 0.25 234.305 ;
			LAYER	M3 ;
			RECT	0 234.205 0.25 234.305 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[65]

	PIN WENB[66]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 237.085 0.25 237.185 ;
			LAYER	M2 ;
			RECT	0 237.085 0.25 237.185 ;
			LAYER	M3 ;
			RECT	0 237.085 0.25 237.185 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[66]

	PIN WENB[67]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 239.965 0.25 240.065 ;
			LAYER	M2 ;
			RECT	0 239.965 0.25 240.065 ;
			LAYER	M3 ;
			RECT	0 239.965 0.25 240.065 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[67]

	PIN WENB[68]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 242.845 0.25 242.945 ;
			LAYER	M2 ;
			RECT	0 242.845 0.25 242.945 ;
			LAYER	M3 ;
			RECT	0 242.845 0.25 242.945 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[68]

	PIN WENB[69]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 245.725 0.25 245.825 ;
			LAYER	M2 ;
			RECT	0 245.725 0.25 245.825 ;
			LAYER	M3 ;
			RECT	0 245.725 0.25 245.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[69]

	PIN WENB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 19.275 0.25 19.375 ;
			LAYER	M2 ;
			RECT	0 19.275 0.25 19.375 ;
			LAYER	M3 ;
			RECT	0 19.275 0.25 19.375 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[6]

	PIN WENB[70]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 248.605 0.25 248.705 ;
			LAYER	M2 ;
			RECT	0 248.605 0.25 248.705 ;
			LAYER	M3 ;
			RECT	0 248.605 0.25 248.705 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[70]

	PIN WENB[71]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 251.485 0.25 251.585 ;
			LAYER	M2 ;
			RECT	0 251.485 0.25 251.585 ;
			LAYER	M3 ;
			RECT	0 251.485 0.25 251.585 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[71]

	PIN WENB[72]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 254.365 0.25 254.465 ;
			LAYER	M2 ;
			RECT	0 254.365 0.25 254.465 ;
			LAYER	M3 ;
			RECT	0 254.365 0.25 254.465 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[72]

	PIN WENB[73]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 257.245 0.25 257.345 ;
			LAYER	M2 ;
			RECT	0 257.245 0.25 257.345 ;
			LAYER	M3 ;
			RECT	0 257.245 0.25 257.345 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[73]

	PIN WENB[74]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 260.125 0.25 260.225 ;
			LAYER	M2 ;
			RECT	0 260.125 0.25 260.225 ;
			LAYER	M3 ;
			RECT	0 260.125 0.25 260.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[74]

	PIN WENB[75]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 263.005 0.25 263.105 ;
			LAYER	M2 ;
			RECT	0 263.005 0.25 263.105 ;
			LAYER	M3 ;
			RECT	0 263.005 0.25 263.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[75]

	PIN WENB[76]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 265.885 0.25 265.985 ;
			LAYER	M2 ;
			RECT	0 265.885 0.25 265.985 ;
			LAYER	M3 ;
			RECT	0 265.885 0.25 265.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[76]

	PIN WENB[77]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 268.765 0.25 268.865 ;
			LAYER	M2 ;
			RECT	0 268.765 0.25 268.865 ;
			LAYER	M3 ;
			RECT	0 268.765 0.25 268.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[77]

	PIN WENB[78]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 271.645 0.25 271.745 ;
			LAYER	M2 ;
			RECT	0 271.645 0.25 271.745 ;
			LAYER	M3 ;
			RECT	0 271.645 0.25 271.745 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[78]

	PIN WENB[79]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 274.525 0.25 274.625 ;
			LAYER	M2 ;
			RECT	0 274.525 0.25 274.625 ;
			LAYER	M3 ;
			RECT	0 274.525 0.25 274.625 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[79]

	PIN WENB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 22.155 0.25 22.255 ;
			LAYER	M2 ;
			RECT	0 22.155 0.25 22.255 ;
			LAYER	M3 ;
			RECT	0 22.155 0.25 22.255 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[7]

	PIN WENB[80]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 277.405 0.25 277.505 ;
			LAYER	M2 ;
			RECT	0 277.405 0.25 277.505 ;
			LAYER	M3 ;
			RECT	0 277.405 0.25 277.505 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[80]

	PIN WENB[81]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 280.285 0.25 280.385 ;
			LAYER	M2 ;
			RECT	0 280.285 0.25 280.385 ;
			LAYER	M3 ;
			RECT	0 280.285 0.25 280.385 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[81]

	PIN WENB[82]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 283.165 0.25 283.265 ;
			LAYER	M2 ;
			RECT	0 283.165 0.25 283.265 ;
			LAYER	M3 ;
			RECT	0 283.165 0.25 283.265 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[82]

	PIN WENB[83]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 286.045 0.25 286.145 ;
			LAYER	M2 ;
			RECT	0 286.045 0.25 286.145 ;
			LAYER	M3 ;
			RECT	0 286.045 0.25 286.145 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[83]

	PIN WENB[84]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 288.925 0.25 289.025 ;
			LAYER	M2 ;
			RECT	0 288.925 0.25 289.025 ;
			LAYER	M3 ;
			RECT	0 288.925 0.25 289.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[84]

	PIN WENB[85]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 291.805 0.25 291.905 ;
			LAYER	M2 ;
			RECT	0 291.805 0.25 291.905 ;
			LAYER	M3 ;
			RECT	0 291.805 0.25 291.905 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[85]

	PIN WENB[86]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 294.685 0.25 294.785 ;
			LAYER	M2 ;
			RECT	0 294.685 0.25 294.785 ;
			LAYER	M3 ;
			RECT	0 294.685 0.25 294.785 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[86]

	PIN WENB[87]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 297.565 0.25 297.665 ;
			LAYER	M2 ;
			RECT	0 297.565 0.25 297.665 ;
			LAYER	M3 ;
			RECT	0 297.565 0.25 297.665 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[87]

	PIN WENB[88]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 300.445 0.25 300.545 ;
			LAYER	M2 ;
			RECT	0 300.445 0.25 300.545 ;
			LAYER	M3 ;
			RECT	0 300.445 0.25 300.545 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[88]

	PIN WENB[89]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 303.325 0.25 303.425 ;
			LAYER	M2 ;
			RECT	0 303.325 0.25 303.425 ;
			LAYER	M3 ;
			RECT	0 303.325 0.25 303.425 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[89]

	PIN WENB[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 25.035 0.25 25.135 ;
			LAYER	M2 ;
			RECT	0 25.035 0.25 25.135 ;
			LAYER	M3 ;
			RECT	0 25.035 0.25 25.135 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[8]

	PIN WENB[90]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 306.205 0.25 306.305 ;
			LAYER	M2 ;
			RECT	0 306.205 0.25 306.305 ;
			LAYER	M3 ;
			RECT	0 306.205 0.25 306.305 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[90]

	PIN WENB[91]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 309.085 0.25 309.185 ;
			LAYER	M2 ;
			RECT	0 309.085 0.25 309.185 ;
			LAYER	M3 ;
			RECT	0 309.085 0.25 309.185 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[91]

	PIN WENB[92]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 311.965 0.25 312.065 ;
			LAYER	M2 ;
			RECT	0 311.965 0.25 312.065 ;
			LAYER	M3 ;
			RECT	0 311.965 0.25 312.065 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[92]

	PIN WENB[93]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 314.845 0.25 314.945 ;
			LAYER	M2 ;
			RECT	0 314.845 0.25 314.945 ;
			LAYER	M3 ;
			RECT	0 314.845 0.25 314.945 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[93]

	PIN WENB[94]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 317.725 0.25 317.825 ;
			LAYER	M2 ;
			RECT	0 317.725 0.25 317.825 ;
			LAYER	M3 ;
			RECT	0 317.725 0.25 317.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[94]

	PIN WENB[95]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 320.605 0.25 320.705 ;
			LAYER	M2 ;
			RECT	0 320.605 0.25 320.705 ;
			LAYER	M3 ;
			RECT	0 320.605 0.25 320.705 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[95]

	PIN WENB[96]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 323.485 0.25 323.585 ;
			LAYER	M2 ;
			RECT	0 323.485 0.25 323.585 ;
			LAYER	M3 ;
			RECT	0 323.485 0.25 323.585 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[96]

	PIN WENB[97]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 326.365 0.25 326.465 ;
			LAYER	M2 ;
			RECT	0 326.365 0.25 326.465 ;
			LAYER	M3 ;
			RECT	0 326.365 0.25 326.465 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[97]

	PIN WENB[98]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 329.245 0.25 329.345 ;
			LAYER	M2 ;
			RECT	0 329.245 0.25 329.345 ;
			LAYER	M3 ;
			RECT	0 329.245 0.25 329.345 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[98]

	PIN WENB[99]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 332.125 0.25 332.225 ;
			LAYER	M2 ;
			RECT	0 332.125 0.25 332.225 ;
			LAYER	M3 ;
			RECT	0 332.125 0.25 332.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[99]

	PIN WENB[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 27.915 0.25 28.015 ;
			LAYER	M2 ;
			RECT	0 27.915 0.25 28.015 ;
			LAYER	M3 ;
			RECT	0 27.915 0.25 28.015 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENB[9]

	PIN WENYB[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 1.73 0.25 1.83 ;
			LAYER	M2 ;
			RECT	0 1.73 0.25 1.83 ;
			LAYER	M3 ;
			RECT	0 1.73 0.25 1.83 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[0]

	PIN WENYB[100]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 335.27 0.25 335.37 ;
			LAYER	M2 ;
			RECT	0 335.27 0.25 335.37 ;
			LAYER	M3 ;
			RECT	0 335.27 0.25 335.37 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[100]

	PIN WENYB[101]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 338.15 0.25 338.25 ;
			LAYER	M2 ;
			RECT	0 338.15 0.25 338.25 ;
			LAYER	M3 ;
			RECT	0 338.15 0.25 338.25 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[101]

	PIN WENYB[102]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 341.03 0.25 341.13 ;
			LAYER	M2 ;
			RECT	0 341.03 0.25 341.13 ;
			LAYER	M3 ;
			RECT	0 341.03 0.25 341.13 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[102]

	PIN WENYB[103]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 343.91 0.25 344.01 ;
			LAYER	M2 ;
			RECT	0 343.91 0.25 344.01 ;
			LAYER	M3 ;
			RECT	0 343.91 0.25 344.01 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[103]

	PIN WENYB[104]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 346.79 0.25 346.89 ;
			LAYER	M2 ;
			RECT	0 346.79 0.25 346.89 ;
			LAYER	M3 ;
			RECT	0 346.79 0.25 346.89 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[104]

	PIN WENYB[105]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 349.67 0.25 349.77 ;
			LAYER	M2 ;
			RECT	0 349.67 0.25 349.77 ;
			LAYER	M3 ;
			RECT	0 349.67 0.25 349.77 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[105]

	PIN WENYB[106]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 352.55 0.25 352.65 ;
			LAYER	M2 ;
			RECT	0 352.55 0.25 352.65 ;
			LAYER	M3 ;
			RECT	0 352.55 0.25 352.65 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[106]

	PIN WENYB[107]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 355.43 0.25 355.53 ;
			LAYER	M2 ;
			RECT	0 355.43 0.25 355.53 ;
			LAYER	M3 ;
			RECT	0 355.43 0.25 355.53 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[107]

	PIN WENYB[108]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 358.31 0.25 358.41 ;
			LAYER	M2 ;
			RECT	0 358.31 0.25 358.41 ;
			LAYER	M3 ;
			RECT	0 358.31 0.25 358.41 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[108]

	PIN WENYB[109]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 361.19 0.25 361.29 ;
			LAYER	M2 ;
			RECT	0 361.19 0.25 361.29 ;
			LAYER	M3 ;
			RECT	0 361.19 0.25 361.29 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[109]

	PIN WENYB[10]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 30.53 0.25 30.63 ;
			LAYER	M2 ;
			RECT	0 30.53 0.25 30.63 ;
			LAYER	M3 ;
			RECT	0 30.53 0.25 30.63 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[10]

	PIN WENYB[110]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 364.07 0.25 364.17 ;
			LAYER	M2 ;
			RECT	0 364.07 0.25 364.17 ;
			LAYER	M3 ;
			RECT	0 364.07 0.25 364.17 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[110]

	PIN WENYB[111]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 366.95 0.25 367.05 ;
			LAYER	M2 ;
			RECT	0 366.95 0.25 367.05 ;
			LAYER	M3 ;
			RECT	0 366.95 0.25 367.05 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[111]

	PIN WENYB[112]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 369.83 0.25 369.93 ;
			LAYER	M2 ;
			RECT	0 369.83 0.25 369.93 ;
			LAYER	M3 ;
			RECT	0 369.83 0.25 369.93 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[112]

	PIN WENYB[113]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 372.71 0.25 372.81 ;
			LAYER	M2 ;
			RECT	0 372.71 0.25 372.81 ;
			LAYER	M3 ;
			RECT	0 372.71 0.25 372.81 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[113]

	PIN WENYB[114]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 375.59 0.25 375.69 ;
			LAYER	M2 ;
			RECT	0 375.59 0.25 375.69 ;
			LAYER	M3 ;
			RECT	0 375.59 0.25 375.69 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[114]

	PIN WENYB[115]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 378.47 0.25 378.57 ;
			LAYER	M2 ;
			RECT	0 378.47 0.25 378.57 ;
			LAYER	M3 ;
			RECT	0 378.47 0.25 378.57 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[115]

	PIN WENYB[116]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 381.35 0.25 381.45 ;
			LAYER	M2 ;
			RECT	0 381.35 0.25 381.45 ;
			LAYER	M3 ;
			RECT	0 381.35 0.25 381.45 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[116]

	PIN WENYB[117]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 384.23 0.25 384.33 ;
			LAYER	M2 ;
			RECT	0 384.23 0.25 384.33 ;
			LAYER	M3 ;
			RECT	0 384.23 0.25 384.33 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[117]

	PIN WENYB[118]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 387.11 0.25 387.21 ;
			LAYER	M2 ;
			RECT	0 387.11 0.25 387.21 ;
			LAYER	M3 ;
			RECT	0 387.11 0.25 387.21 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[118]

	PIN WENYB[119]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 389.99 0.25 390.09 ;
			LAYER	M2 ;
			RECT	0 389.99 0.25 390.09 ;
			LAYER	M3 ;
			RECT	0 389.99 0.25 390.09 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[119]

	PIN WENYB[11]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 33.41 0.25 33.51 ;
			LAYER	M2 ;
			RECT	0 33.41 0.25 33.51 ;
			LAYER	M3 ;
			RECT	0 33.41 0.25 33.51 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[11]

	PIN WENYB[120]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 392.87 0.25 392.97 ;
			LAYER	M2 ;
			RECT	0 392.87 0.25 392.97 ;
			LAYER	M3 ;
			RECT	0 392.87 0.25 392.97 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[120]

	PIN WENYB[121]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 395.75 0.25 395.85 ;
			LAYER	M2 ;
			RECT	0 395.75 0.25 395.85 ;
			LAYER	M3 ;
			RECT	0 395.75 0.25 395.85 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[121]

	PIN WENYB[122]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 398.63 0.25 398.73 ;
			LAYER	M2 ;
			RECT	0 398.63 0.25 398.73 ;
			LAYER	M3 ;
			RECT	0 398.63 0.25 398.73 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[122]

	PIN WENYB[123]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 401.51 0.25 401.61 ;
			LAYER	M2 ;
			RECT	0 401.51 0.25 401.61 ;
			LAYER	M3 ;
			RECT	0 401.51 0.25 401.61 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[123]

	PIN WENYB[124]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 404.39 0.25 404.49 ;
			LAYER	M2 ;
			RECT	0 404.39 0.25 404.49 ;
			LAYER	M3 ;
			RECT	0 404.39 0.25 404.49 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[124]

	PIN WENYB[125]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 407.27 0.25 407.37 ;
			LAYER	M2 ;
			RECT	0 407.27 0.25 407.37 ;
			LAYER	M3 ;
			RECT	0 407.27 0.25 407.37 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[125]

	PIN WENYB[126]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 410.15 0.25 410.25 ;
			LAYER	M2 ;
			RECT	0 410.15 0.25 410.25 ;
			LAYER	M3 ;
			RECT	0 410.15 0.25 410.25 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[126]

	PIN WENYB[127]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 413.03 0.25 413.13 ;
			LAYER	M2 ;
			RECT	0 413.03 0.25 413.13 ;
			LAYER	M3 ;
			RECT	0 413.03 0.25 413.13 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[127]

	PIN WENYB[12]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 36.29 0.25 36.39 ;
			LAYER	M2 ;
			RECT	0 36.29 0.25 36.39 ;
			LAYER	M3 ;
			RECT	0 36.29 0.25 36.39 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[12]

	PIN WENYB[13]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 39.17 0.25 39.27 ;
			LAYER	M2 ;
			RECT	0 39.17 0.25 39.27 ;
			LAYER	M3 ;
			RECT	0 39.17 0.25 39.27 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[13]

	PIN WENYB[14]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 42.05 0.25 42.15 ;
			LAYER	M2 ;
			RECT	0 42.05 0.25 42.15 ;
			LAYER	M3 ;
			RECT	0 42.05 0.25 42.15 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[14]

	PIN WENYB[15]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 44.93 0.25 45.03 ;
			LAYER	M2 ;
			RECT	0 44.93 0.25 45.03 ;
			LAYER	M3 ;
			RECT	0 44.93 0.25 45.03 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[15]

	PIN WENYB[16]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 47.81 0.25 47.91 ;
			LAYER	M2 ;
			RECT	0 47.81 0.25 47.91 ;
			LAYER	M3 ;
			RECT	0 47.81 0.25 47.91 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[16]

	PIN WENYB[17]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 50.69 0.25 50.79 ;
			LAYER	M2 ;
			RECT	0 50.69 0.25 50.79 ;
			LAYER	M3 ;
			RECT	0 50.69 0.25 50.79 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[17]

	PIN WENYB[18]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 53.57 0.25 53.67 ;
			LAYER	M2 ;
			RECT	0 53.57 0.25 53.67 ;
			LAYER	M3 ;
			RECT	0 53.57 0.25 53.67 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[18]

	PIN WENYB[19]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 56.45 0.25 56.55 ;
			LAYER	M2 ;
			RECT	0 56.45 0.25 56.55 ;
			LAYER	M3 ;
			RECT	0 56.45 0.25 56.55 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[19]

	PIN WENYB[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 4.61 0.25 4.71 ;
			LAYER	M2 ;
			RECT	0 4.61 0.25 4.71 ;
			LAYER	M3 ;
			RECT	0 4.61 0.25 4.71 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[1]

	PIN WENYB[20]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 59.33 0.25 59.43 ;
			LAYER	M2 ;
			RECT	0 59.33 0.25 59.43 ;
			LAYER	M3 ;
			RECT	0 59.33 0.25 59.43 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[20]

	PIN WENYB[21]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 62.21 0.25 62.31 ;
			LAYER	M2 ;
			RECT	0 62.21 0.25 62.31 ;
			LAYER	M3 ;
			RECT	0 62.21 0.25 62.31 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[21]

	PIN WENYB[22]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 65.09 0.25 65.19 ;
			LAYER	M2 ;
			RECT	0 65.09 0.25 65.19 ;
			LAYER	M3 ;
			RECT	0 65.09 0.25 65.19 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[22]

	PIN WENYB[23]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 67.97 0.25 68.07 ;
			LAYER	M2 ;
			RECT	0 67.97 0.25 68.07 ;
			LAYER	M3 ;
			RECT	0 67.97 0.25 68.07 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[23]

	PIN WENYB[24]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 70.85 0.25 70.95 ;
			LAYER	M2 ;
			RECT	0 70.85 0.25 70.95 ;
			LAYER	M3 ;
			RECT	0 70.85 0.25 70.95 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[24]

	PIN WENYB[25]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 73.73 0.25 73.83 ;
			LAYER	M2 ;
			RECT	0 73.73 0.25 73.83 ;
			LAYER	M3 ;
			RECT	0 73.73 0.25 73.83 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[25]

	PIN WENYB[26]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 76.61 0.25 76.71 ;
			LAYER	M2 ;
			RECT	0 76.61 0.25 76.71 ;
			LAYER	M3 ;
			RECT	0 76.61 0.25 76.71 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[26]

	PIN WENYB[27]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 79.49 0.25 79.59 ;
			LAYER	M2 ;
			RECT	0 79.49 0.25 79.59 ;
			LAYER	M3 ;
			RECT	0 79.49 0.25 79.59 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[27]

	PIN WENYB[28]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 82.37 0.25 82.47 ;
			LAYER	M2 ;
			RECT	0 82.37 0.25 82.47 ;
			LAYER	M3 ;
			RECT	0 82.37 0.25 82.47 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[28]

	PIN WENYB[29]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 85.25 0.25 85.35 ;
			LAYER	M2 ;
			RECT	0 85.25 0.25 85.35 ;
			LAYER	M3 ;
			RECT	0 85.25 0.25 85.35 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[29]

	PIN WENYB[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 7.49 0.25 7.59 ;
			LAYER	M2 ;
			RECT	0 7.49 0.25 7.59 ;
			LAYER	M3 ;
			RECT	0 7.49 0.25 7.59 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[2]

	PIN WENYB[30]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 88.13 0.25 88.23 ;
			LAYER	M2 ;
			RECT	0 88.13 0.25 88.23 ;
			LAYER	M3 ;
			RECT	0 88.13 0.25 88.23 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[30]

	PIN WENYB[31]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 91.01 0.25 91.11 ;
			LAYER	M2 ;
			RECT	0 91.01 0.25 91.11 ;
			LAYER	M3 ;
			RECT	0 91.01 0.25 91.11 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[31]

	PIN WENYB[32]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 93.89 0.25 93.99 ;
			LAYER	M2 ;
			RECT	0 93.89 0.25 93.99 ;
			LAYER	M3 ;
			RECT	0 93.89 0.25 93.99 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[32]

	PIN WENYB[33]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 96.77 0.25 96.87 ;
			LAYER	M2 ;
			RECT	0 96.77 0.25 96.87 ;
			LAYER	M3 ;
			RECT	0 96.77 0.25 96.87 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[33]

	PIN WENYB[34]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 99.65 0.25 99.75 ;
			LAYER	M2 ;
			RECT	0 99.65 0.25 99.75 ;
			LAYER	M3 ;
			RECT	0 99.65 0.25 99.75 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[34]

	PIN WENYB[35]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 102.53 0.25 102.63 ;
			LAYER	M2 ;
			RECT	0 102.53 0.25 102.63 ;
			LAYER	M3 ;
			RECT	0 102.53 0.25 102.63 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[35]

	PIN WENYB[36]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 105.41 0.25 105.51 ;
			LAYER	M2 ;
			RECT	0 105.41 0.25 105.51 ;
			LAYER	M3 ;
			RECT	0 105.41 0.25 105.51 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[36]

	PIN WENYB[37]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 108.29 0.25 108.39 ;
			LAYER	M2 ;
			RECT	0 108.29 0.25 108.39 ;
			LAYER	M3 ;
			RECT	0 108.29 0.25 108.39 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[37]

	PIN WENYB[38]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 111.17 0.25 111.27 ;
			LAYER	M2 ;
			RECT	0 111.17 0.25 111.27 ;
			LAYER	M3 ;
			RECT	0 111.17 0.25 111.27 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[38]

	PIN WENYB[39]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 114.05 0.25 114.15 ;
			LAYER	M2 ;
			RECT	0 114.05 0.25 114.15 ;
			LAYER	M3 ;
			RECT	0 114.05 0.25 114.15 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[39]

	PIN WENYB[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 10.37 0.25 10.47 ;
			LAYER	M2 ;
			RECT	0 10.37 0.25 10.47 ;
			LAYER	M3 ;
			RECT	0 10.37 0.25 10.47 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[3]

	PIN WENYB[40]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 116.93 0.25 117.03 ;
			LAYER	M2 ;
			RECT	0 116.93 0.25 117.03 ;
			LAYER	M3 ;
			RECT	0 116.93 0.25 117.03 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[40]

	PIN WENYB[41]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 119.81 0.25 119.91 ;
			LAYER	M2 ;
			RECT	0 119.81 0.25 119.91 ;
			LAYER	M3 ;
			RECT	0 119.81 0.25 119.91 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[41]

	PIN WENYB[42]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 122.69 0.25 122.79 ;
			LAYER	M2 ;
			RECT	0 122.69 0.25 122.79 ;
			LAYER	M3 ;
			RECT	0 122.69 0.25 122.79 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[42]

	PIN WENYB[43]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 125.57 0.25 125.67 ;
			LAYER	M2 ;
			RECT	0 125.57 0.25 125.67 ;
			LAYER	M3 ;
			RECT	0 125.57 0.25 125.67 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[43]

	PIN WENYB[44]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 128.45 0.25 128.55 ;
			LAYER	M2 ;
			RECT	0 128.45 0.25 128.55 ;
			LAYER	M3 ;
			RECT	0 128.45 0.25 128.55 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[44]

	PIN WENYB[45]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 131.33 0.25 131.43 ;
			LAYER	M2 ;
			RECT	0 131.33 0.25 131.43 ;
			LAYER	M3 ;
			RECT	0 131.33 0.25 131.43 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[45]

	PIN WENYB[46]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 134.21 0.25 134.31 ;
			LAYER	M2 ;
			RECT	0 134.21 0.25 134.31 ;
			LAYER	M3 ;
			RECT	0 134.21 0.25 134.31 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[46]

	PIN WENYB[47]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 137.09 0.25 137.19 ;
			LAYER	M2 ;
			RECT	0 137.09 0.25 137.19 ;
			LAYER	M3 ;
			RECT	0 137.09 0.25 137.19 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[47]

	PIN WENYB[48]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 139.97 0.25 140.07 ;
			LAYER	M2 ;
			RECT	0 139.97 0.25 140.07 ;
			LAYER	M3 ;
			RECT	0 139.97 0.25 140.07 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[48]

	PIN WENYB[49]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 142.85 0.25 142.95 ;
			LAYER	M2 ;
			RECT	0 142.85 0.25 142.95 ;
			LAYER	M3 ;
			RECT	0 142.85 0.25 142.95 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[49]

	PIN WENYB[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 13.25 0.25 13.35 ;
			LAYER	M2 ;
			RECT	0 13.25 0.25 13.35 ;
			LAYER	M3 ;
			RECT	0 13.25 0.25 13.35 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[4]

	PIN WENYB[50]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 145.73 0.25 145.83 ;
			LAYER	M2 ;
			RECT	0 145.73 0.25 145.83 ;
			LAYER	M3 ;
			RECT	0 145.73 0.25 145.83 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[50]

	PIN WENYB[51]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 148.61 0.25 148.71 ;
			LAYER	M2 ;
			RECT	0 148.61 0.25 148.71 ;
			LAYER	M3 ;
			RECT	0 148.61 0.25 148.71 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[51]

	PIN WENYB[52]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 151.49 0.25 151.59 ;
			LAYER	M2 ;
			RECT	0 151.49 0.25 151.59 ;
			LAYER	M3 ;
			RECT	0 151.49 0.25 151.59 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[52]

	PIN WENYB[53]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 154.37 0.25 154.47 ;
			LAYER	M2 ;
			RECT	0 154.37 0.25 154.47 ;
			LAYER	M3 ;
			RECT	0 154.37 0.25 154.47 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[53]

	PIN WENYB[54]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 157.25 0.25 157.35 ;
			LAYER	M2 ;
			RECT	0 157.25 0.25 157.35 ;
			LAYER	M3 ;
			RECT	0 157.25 0.25 157.35 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[54]

	PIN WENYB[55]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 160.13 0.25 160.23 ;
			LAYER	M2 ;
			RECT	0 160.13 0.25 160.23 ;
			LAYER	M3 ;
			RECT	0 160.13 0.25 160.23 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[55]

	PIN WENYB[56]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 163.01 0.25 163.11 ;
			LAYER	M2 ;
			RECT	0 163.01 0.25 163.11 ;
			LAYER	M3 ;
			RECT	0 163.01 0.25 163.11 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[56]

	PIN WENYB[57]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 165.89 0.25 165.99 ;
			LAYER	M2 ;
			RECT	0 165.89 0.25 165.99 ;
			LAYER	M3 ;
			RECT	0 165.89 0.25 165.99 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[57]

	PIN WENYB[58]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 168.77 0.25 168.87 ;
			LAYER	M2 ;
			RECT	0 168.77 0.25 168.87 ;
			LAYER	M3 ;
			RECT	0 168.77 0.25 168.87 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[58]

	PIN WENYB[59]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 171.65 0.25 171.75 ;
			LAYER	M2 ;
			RECT	0 171.65 0.25 171.75 ;
			LAYER	M3 ;
			RECT	0 171.65 0.25 171.75 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[59]

	PIN WENYB[5]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 16.13 0.25 16.23 ;
			LAYER	M2 ;
			RECT	0 16.13 0.25 16.23 ;
			LAYER	M3 ;
			RECT	0 16.13 0.25 16.23 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[5]

	PIN WENYB[60]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 174.53 0.25 174.63 ;
			LAYER	M2 ;
			RECT	0 174.53 0.25 174.63 ;
			LAYER	M3 ;
			RECT	0 174.53 0.25 174.63 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[60]

	PIN WENYB[61]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 177.41 0.25 177.51 ;
			LAYER	M2 ;
			RECT	0 177.41 0.25 177.51 ;
			LAYER	M3 ;
			RECT	0 177.41 0.25 177.51 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[61]

	PIN WENYB[62]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 180.29 0.25 180.39 ;
			LAYER	M2 ;
			RECT	0 180.29 0.25 180.39 ;
			LAYER	M3 ;
			RECT	0 180.29 0.25 180.39 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[62]

	PIN WENYB[63]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 183.17 0.25 183.27 ;
			LAYER	M2 ;
			RECT	0 183.17 0.25 183.27 ;
			LAYER	M3 ;
			RECT	0 183.17 0.25 183.27 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[63]

	PIN WENYB[64]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 231.59 0.25 231.69 ;
			LAYER	M2 ;
			RECT	0 231.59 0.25 231.69 ;
			LAYER	M3 ;
			RECT	0 231.59 0.25 231.69 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[64]

	PIN WENYB[65]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 234.47 0.25 234.57 ;
			LAYER	M2 ;
			RECT	0 234.47 0.25 234.57 ;
			LAYER	M3 ;
			RECT	0 234.47 0.25 234.57 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[65]

	PIN WENYB[66]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 237.35 0.25 237.45 ;
			LAYER	M2 ;
			RECT	0 237.35 0.25 237.45 ;
			LAYER	M3 ;
			RECT	0 237.35 0.25 237.45 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[66]

	PIN WENYB[67]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 240.23 0.25 240.33 ;
			LAYER	M2 ;
			RECT	0 240.23 0.25 240.33 ;
			LAYER	M3 ;
			RECT	0 240.23 0.25 240.33 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[67]

	PIN WENYB[68]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 243.11 0.25 243.21 ;
			LAYER	M2 ;
			RECT	0 243.11 0.25 243.21 ;
			LAYER	M3 ;
			RECT	0 243.11 0.25 243.21 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[68]

	PIN WENYB[69]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 245.99 0.25 246.09 ;
			LAYER	M2 ;
			RECT	0 245.99 0.25 246.09 ;
			LAYER	M3 ;
			RECT	0 245.99 0.25 246.09 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[69]

	PIN WENYB[6]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 19.01 0.25 19.11 ;
			LAYER	M2 ;
			RECT	0 19.01 0.25 19.11 ;
			LAYER	M3 ;
			RECT	0 19.01 0.25 19.11 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[6]

	PIN WENYB[70]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 248.87 0.25 248.97 ;
			LAYER	M2 ;
			RECT	0 248.87 0.25 248.97 ;
			LAYER	M3 ;
			RECT	0 248.87 0.25 248.97 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[70]

	PIN WENYB[71]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 251.75 0.25 251.85 ;
			LAYER	M2 ;
			RECT	0 251.75 0.25 251.85 ;
			LAYER	M3 ;
			RECT	0 251.75 0.25 251.85 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[71]

	PIN WENYB[72]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 254.63 0.25 254.73 ;
			LAYER	M2 ;
			RECT	0 254.63 0.25 254.73 ;
			LAYER	M3 ;
			RECT	0 254.63 0.25 254.73 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[72]

	PIN WENYB[73]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 257.51 0.25 257.61 ;
			LAYER	M2 ;
			RECT	0 257.51 0.25 257.61 ;
			LAYER	M3 ;
			RECT	0 257.51 0.25 257.61 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[73]

	PIN WENYB[74]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 260.39 0.25 260.49 ;
			LAYER	M2 ;
			RECT	0 260.39 0.25 260.49 ;
			LAYER	M3 ;
			RECT	0 260.39 0.25 260.49 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[74]

	PIN WENYB[75]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 263.27 0.25 263.37 ;
			LAYER	M2 ;
			RECT	0 263.27 0.25 263.37 ;
			LAYER	M3 ;
			RECT	0 263.27 0.25 263.37 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[75]

	PIN WENYB[76]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 266.15 0.25 266.25 ;
			LAYER	M2 ;
			RECT	0 266.15 0.25 266.25 ;
			LAYER	M3 ;
			RECT	0 266.15 0.25 266.25 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[76]

	PIN WENYB[77]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 269.03 0.25 269.13 ;
			LAYER	M2 ;
			RECT	0 269.03 0.25 269.13 ;
			LAYER	M3 ;
			RECT	0 269.03 0.25 269.13 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[77]

	PIN WENYB[78]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 271.91 0.25 272.01 ;
			LAYER	M2 ;
			RECT	0 271.91 0.25 272.01 ;
			LAYER	M3 ;
			RECT	0 271.91 0.25 272.01 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[78]

	PIN WENYB[79]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 274.79 0.25 274.89 ;
			LAYER	M2 ;
			RECT	0 274.79 0.25 274.89 ;
			LAYER	M3 ;
			RECT	0 274.79 0.25 274.89 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[79]

	PIN WENYB[7]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 21.89 0.25 21.99 ;
			LAYER	M2 ;
			RECT	0 21.89 0.25 21.99 ;
			LAYER	M3 ;
			RECT	0 21.89 0.25 21.99 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[7]

	PIN WENYB[80]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 277.67 0.25 277.77 ;
			LAYER	M2 ;
			RECT	0 277.67 0.25 277.77 ;
			LAYER	M3 ;
			RECT	0 277.67 0.25 277.77 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[80]

	PIN WENYB[81]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 280.55 0.25 280.65 ;
			LAYER	M2 ;
			RECT	0 280.55 0.25 280.65 ;
			LAYER	M3 ;
			RECT	0 280.55 0.25 280.65 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[81]

	PIN WENYB[82]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 283.43 0.25 283.53 ;
			LAYER	M2 ;
			RECT	0 283.43 0.25 283.53 ;
			LAYER	M3 ;
			RECT	0 283.43 0.25 283.53 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[82]

	PIN WENYB[83]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 286.31 0.25 286.41 ;
			LAYER	M2 ;
			RECT	0 286.31 0.25 286.41 ;
			LAYER	M3 ;
			RECT	0 286.31 0.25 286.41 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[83]

	PIN WENYB[84]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 289.19 0.25 289.29 ;
			LAYER	M2 ;
			RECT	0 289.19 0.25 289.29 ;
			LAYER	M3 ;
			RECT	0 289.19 0.25 289.29 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[84]

	PIN WENYB[85]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 292.07 0.25 292.17 ;
			LAYER	M2 ;
			RECT	0 292.07 0.25 292.17 ;
			LAYER	M3 ;
			RECT	0 292.07 0.25 292.17 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[85]

	PIN WENYB[86]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 294.95 0.25 295.05 ;
			LAYER	M2 ;
			RECT	0 294.95 0.25 295.05 ;
			LAYER	M3 ;
			RECT	0 294.95 0.25 295.05 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[86]

	PIN WENYB[87]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 297.83 0.25 297.93 ;
			LAYER	M2 ;
			RECT	0 297.83 0.25 297.93 ;
			LAYER	M3 ;
			RECT	0 297.83 0.25 297.93 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[87]

	PIN WENYB[88]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 300.71 0.25 300.81 ;
			LAYER	M2 ;
			RECT	0 300.71 0.25 300.81 ;
			LAYER	M3 ;
			RECT	0 300.71 0.25 300.81 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[88]

	PIN WENYB[89]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 303.59 0.25 303.69 ;
			LAYER	M2 ;
			RECT	0 303.59 0.25 303.69 ;
			LAYER	M3 ;
			RECT	0 303.59 0.25 303.69 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[89]

	PIN WENYB[8]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 24.77 0.25 24.87 ;
			LAYER	M2 ;
			RECT	0 24.77 0.25 24.87 ;
			LAYER	M3 ;
			RECT	0 24.77 0.25 24.87 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[8]

	PIN WENYB[90]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 306.47 0.25 306.57 ;
			LAYER	M2 ;
			RECT	0 306.47 0.25 306.57 ;
			LAYER	M3 ;
			RECT	0 306.47 0.25 306.57 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[90]

	PIN WENYB[91]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 309.35 0.25 309.45 ;
			LAYER	M2 ;
			RECT	0 309.35 0.25 309.45 ;
			LAYER	M3 ;
			RECT	0 309.35 0.25 309.45 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[91]

	PIN WENYB[92]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 312.23 0.25 312.33 ;
			LAYER	M2 ;
			RECT	0 312.23 0.25 312.33 ;
			LAYER	M3 ;
			RECT	0 312.23 0.25 312.33 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[92]

	PIN WENYB[93]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 315.11 0.25 315.21 ;
			LAYER	M2 ;
			RECT	0 315.11 0.25 315.21 ;
			LAYER	M3 ;
			RECT	0 315.11 0.25 315.21 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[93]

	PIN WENYB[94]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 317.99 0.25 318.09 ;
			LAYER	M2 ;
			RECT	0 317.99 0.25 318.09 ;
			LAYER	M3 ;
			RECT	0 317.99 0.25 318.09 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[94]

	PIN WENYB[95]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 320.87 0.25 320.97 ;
			LAYER	M2 ;
			RECT	0 320.87 0.25 320.97 ;
			LAYER	M3 ;
			RECT	0 320.87 0.25 320.97 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[95]

	PIN WENYB[96]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 323.75 0.25 323.85 ;
			LAYER	M2 ;
			RECT	0 323.75 0.25 323.85 ;
			LAYER	M3 ;
			RECT	0 323.75 0.25 323.85 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[96]

	PIN WENYB[97]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 326.63 0.25 326.73 ;
			LAYER	M2 ;
			RECT	0 326.63 0.25 326.73 ;
			LAYER	M3 ;
			RECT	0 326.63 0.25 326.73 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[97]

	PIN WENYB[98]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 329.51 0.25 329.61 ;
			LAYER	M2 ;
			RECT	0 329.51 0.25 329.61 ;
			LAYER	M3 ;
			RECT	0 329.51 0.25 329.61 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[98]

	PIN WENYB[99]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 332.39 0.25 332.49 ;
			LAYER	M2 ;
			RECT	0 332.39 0.25 332.49 ;
			LAYER	M3 ;
			RECT	0 332.39 0.25 332.49 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[99]

	PIN WENYB[9]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 27.65 0.25 27.75 ;
			LAYER	M2 ;
			RECT	0 27.65 0.25 27.75 ;
			LAYER	M3 ;
			RECT	0 27.65 0.25 27.75 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END WENYB[9]

	OBS
		LAYER	M1 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0.35 21.655 414.51 ;
		RECT	0 0.56 0.32 1.365 ;
		RECT	0 2.655 0.32 3.16 ;
		RECT	0 3.46 0.32 4.245 ;
		RECT	0 5.535 0.32 6.04 ;
		RECT	0 6.34 0.32 7.125 ;
		RECT	0 8.415 0.32 8.92 ;
		RECT	0 9.22 0.32 10.005 ;
		RECT	0 11.295 0.32 11.8 ;
		RECT	0 12.1 0.32 12.885 ;
		RECT	0 14.175 0.32 14.68 ;
		RECT	0 14.98 0.32 15.765 ;
		RECT	0 17.055 0.32 17.56 ;
		RECT	0 17.86 0.32 18.645 ;
		RECT	0 19.935 0.32 20.44 ;
		RECT	0 20.74 0.32 21.525 ;
		RECT	0 22.815 0.32 23.32 ;
		RECT	0 23.62 0.32 24.405 ;
		RECT	0 25.695 0.32 26.2 ;
		RECT	0 26.5 0.32 27.285 ;
		RECT	0 28.575 0.32 29.08 ;
		RECT	0 29.38 0.32 30.165 ;
		RECT	0 31.455 0.32 31.96 ;
		RECT	0 32.26 0.32 33.045 ;
		RECT	0 34.335 0.32 34.84 ;
		RECT	0 35.14 0.32 35.925 ;
		RECT	0 37.215 0.32 37.72 ;
		RECT	0 38.02 0.32 38.805 ;
		RECT	0 40.095 0.32 40.6 ;
		RECT	0 40.9 0.32 41.685 ;
		RECT	0 42.975 0.32 43.48 ;
		RECT	0 43.78 0.32 44.565 ;
		RECT	0 45.855 0.32 46.36 ;
		RECT	0 46.66 0.32 47.445 ;
		RECT	0 48.735 0.32 49.24 ;
		RECT	0 49.54 0.32 50.325 ;
		RECT	0 51.615 0.32 52.12 ;
		RECT	0 52.42 0.32 53.205 ;
		RECT	0 54.495 0.32 55 ;
		RECT	0 55.3 0.32 56.085 ;
		RECT	0 57.375 0.32 57.88 ;
		RECT	0 58.18 0.32 58.965 ;
		RECT	0 60.255 0.32 60.76 ;
		RECT	0 61.06 0.32 61.845 ;
		RECT	0 63.135 0.32 63.64 ;
		RECT	0 63.94 0.32 64.725 ;
		RECT	0 66.015 0.32 66.52 ;
		RECT	0 66.82 0.32 67.605 ;
		RECT	0 68.895 0.32 69.4 ;
		RECT	0 69.7 0.32 70.485 ;
		RECT	0 71.775 0.32 72.28 ;
		RECT	0 72.58 0.32 73.365 ;
		RECT	0 74.655 0.32 75.16 ;
		RECT	0 75.46 0.32 76.245 ;
		RECT	0 77.535 0.32 78.04 ;
		RECT	0 78.34 0.32 79.125 ;
		RECT	0 80.415 0.32 80.92 ;
		RECT	0 81.22 0.32 82.005 ;
		RECT	0 83.295 0.32 83.8 ;
		RECT	0 84.1 0.32 84.885 ;
		RECT	0 86.175 0.32 86.68 ;
		RECT	0 86.98 0.32 87.765 ;
		RECT	0 89.055 0.32 89.56 ;
		RECT	0 89.86 0.32 90.645 ;
		RECT	0 91.935 0.32 92.44 ;
		RECT	0 92.74 0.32 93.525 ;
		RECT	0 94.815 0.32 95.32 ;
		RECT	0 95.62 0.32 96.405 ;
		RECT	0 97.695 0.32 98.2 ;
		RECT	0 98.5 0.32 99.285 ;
		RECT	0 100.575 0.32 101.08 ;
		RECT	0 101.38 0.32 102.165 ;
		RECT	0 103.455 0.32 103.96 ;
		RECT	0 104.26 0.32 105.045 ;
		RECT	0 106.335 0.32 106.84 ;
		RECT	0 107.14 0.32 107.925 ;
		RECT	0 109.215 0.32 109.72 ;
		RECT	0 110.02 0.32 110.805 ;
		RECT	0 112.095 0.32 112.6 ;
		RECT	0 112.9 0.32 113.685 ;
		RECT	0 114.975 0.32 115.48 ;
		RECT	0 115.78 0.32 116.565 ;
		RECT	0 117.855 0.32 118.36 ;
		RECT	0 118.66 0.32 119.445 ;
		RECT	0 120.735 0.32 121.24 ;
		RECT	0 121.54 0.32 122.325 ;
		RECT	0 123.615 0.32 124.12 ;
		RECT	0 124.42 0.32 125.205 ;
		RECT	0 126.495 0.32 127 ;
		RECT	0 127.3 0.32 128.085 ;
		RECT	0 129.375 0.32 129.88 ;
		RECT	0 130.18 0.32 130.965 ;
		RECT	0 132.255 0.32 132.76 ;
		RECT	0 133.06 0.32 133.845 ;
		RECT	0 135.135 0.32 135.64 ;
		RECT	0 135.94 0.32 136.725 ;
		RECT	0 138.015 0.32 138.52 ;
		RECT	0 138.82 0.32 139.605 ;
		RECT	0 140.895 0.32 141.4 ;
		RECT	0 141.7 0.32 142.485 ;
		RECT	0 143.775 0.32 144.28 ;
		RECT	0 144.58 0.32 145.365 ;
		RECT	0 146.655 0.32 147.16 ;
		RECT	0 147.46 0.32 148.245 ;
		RECT	0 149.535 0.32 150.04 ;
		RECT	0 150.34 0.32 151.125 ;
		RECT	0 152.415 0.32 152.92 ;
		RECT	0 153.22 0.32 154.005 ;
		RECT	0 155.295 0.32 155.8 ;
		RECT	0 156.1 0.32 156.885 ;
		RECT	0 158.175 0.32 158.68 ;
		RECT	0 158.98 0.32 159.765 ;
		RECT	0 161.055 0.32 161.56 ;
		RECT	0 161.86 0.32 162.645 ;
		RECT	0 163.935 0.32 164.44 ;
		RECT	0 164.74 0.32 165.525 ;
		RECT	0 166.815 0.32 167.32 ;
		RECT	0 167.62 0.32 168.405 ;
		RECT	0 169.695 0.32 170.2 ;
		RECT	0 170.5 0.32 171.285 ;
		RECT	0 172.575 0.32 173.08 ;
		RECT	0 173.38 0.32 174.165 ;
		RECT	0 175.455 0.32 175.96 ;
		RECT	0 176.26 0.32 177.045 ;
		RECT	0 178.335 0.32 178.84 ;
		RECT	0 179.14 0.32 179.925 ;
		RECT	0 181.215 0.32 181.72 ;
		RECT	0 182.02 0.32 182.805 ;
		RECT	0 184.095 0.32 184.6 ;
		RECT	0 184.9 0.32 187 ;
		RECT	0 187.3 0.32 187.35 ;
		RECT	0 187.65 0.32 188.01 ;
		RECT	0 188.71 0.32 190.35 ;
		RECT	0 190.955 0.32 191.17 ;
		RECT	0 191.47 0.32 191.575 ;
		RECT	0 191.875 0.32 193.685 ;
		RECT	0 193.985 0.32 194.2 ;
		RECT	0 194.5 0.32 194.605 ;
		RECT	0 194.905 0.32 196.745 ;
		RECT	0 197.045 0.32 197.23 ;
		RECT	0 197.53 0.32 197.635 ;
		RECT	0 197.935 0.32 198.03 ;
		RECT	0 198.33 0.32 198.4 ;
		RECT	0 198.7 0.32 198.775 ;
		RECT	0 199.075 0.32 199.26 ;
		RECT	0 199.97 0.32 201.405 ;
		RECT	0 202.105 0.32 202.29 ;
		RECT	0 202.875 0.32 205.8 ;
		RECT	0 206.5 0.32 206.97 ;
		RECT	0 207.27 0.32 208.635 ;
		RECT	0 208.935 0.32 212.725 ;
		RECT	0 213.26 0.32 213.45 ;
		RECT	0 213.75 0.32 213.825 ;
		RECT	0 214.125 0.32 214.205 ;
		RECT	0 214.505 0.32 215.205 ;
		RECT	0 215.505 0.32 215.995 ;
		RECT	0 216.295 0.32 216.48 ;
		RECT	0 216.78 0.32 216.885 ;
		RECT	0 217.185 0.32 217.65 ;
		RECT	0 217.95 0.32 218.025 ;
		RECT	0 218.325 0.32 218.48 ;
		RECT	0 218.98 0.32 220.225 ;
		RECT	0 220.525 0.32 220.65 ;
		RECT	0 221.16 0.32 221.54 ;
		RECT	0 221.84 0.32 223.68 ;
		RECT	0 223.98 0.32 224.085 ;
		RECT	0 224.385 0.32 224.57 ;
		RECT	0 225.125 0.32 225.6 ;
		RECT	0 225.9 0.32 228.21 ;
		RECT	0 228.51 0.32 228.605 ;
		RECT	0 228.905 0.32 229.15 ;
		RECT	0 229.45 0.32 229.96 ;
		RECT	0 230.26 0.32 230.765 ;
		RECT	0 232.055 0.32 232.84 ;
		RECT	0 233.14 0.32 233.645 ;
		RECT	0 234.935 0.32 235.72 ;
		RECT	0 236.02 0.32 236.525 ;
		RECT	0 237.815 0.32 238.6 ;
		RECT	0 238.9 0.32 239.405 ;
		RECT	0 240.695 0.32 241.48 ;
		RECT	0 241.78 0.32 242.285 ;
		RECT	0 243.575 0.32 244.36 ;
		RECT	0 244.66 0.32 245.165 ;
		RECT	0 246.455 0.32 247.24 ;
		RECT	0 247.54 0.32 248.045 ;
		RECT	0 249.335 0.32 250.12 ;
		RECT	0 250.42 0.32 250.925 ;
		RECT	0 252.215 0.32 253 ;
		RECT	0 253.3 0.32 253.805 ;
		RECT	0 255.095 0.32 255.88 ;
		RECT	0 256.18 0.32 256.685 ;
		RECT	0 257.975 0.32 258.76 ;
		RECT	0 259.06 0.32 259.565 ;
		RECT	0 260.855 0.32 261.64 ;
		RECT	0 261.94 0.32 262.445 ;
		RECT	0 263.735 0.32 264.52 ;
		RECT	0 264.82 0.32 265.325 ;
		RECT	0 266.615 0.32 267.4 ;
		RECT	0 267.7 0.32 268.205 ;
		RECT	0 269.495 0.32 270.28 ;
		RECT	0 270.58 0.32 271.085 ;
		RECT	0 272.375 0.32 273.16 ;
		RECT	0 273.46 0.32 273.965 ;
		RECT	0 275.255 0.32 276.04 ;
		RECT	0 276.34 0.32 276.845 ;
		RECT	0 278.135 0.32 278.92 ;
		RECT	0 279.22 0.32 279.725 ;
		RECT	0 281.015 0.32 281.8 ;
		RECT	0 282.1 0.32 282.605 ;
		RECT	0 283.895 0.32 284.68 ;
		RECT	0 284.98 0.32 285.485 ;
		RECT	0 286.775 0.32 287.56 ;
		RECT	0 287.86 0.32 288.365 ;
		RECT	0 289.655 0.32 290.44 ;
		RECT	0 290.74 0.32 291.245 ;
		RECT	0 292.535 0.32 293.32 ;
		RECT	0 293.62 0.32 294.125 ;
		RECT	0 295.415 0.32 296.2 ;
		RECT	0 296.5 0.32 297.005 ;
		RECT	0 298.295 0.32 299.08 ;
		RECT	0 299.38 0.32 299.885 ;
		RECT	0 301.175 0.32 301.96 ;
		RECT	0 302.26 0.32 302.765 ;
		RECT	0 304.055 0.32 304.84 ;
		RECT	0 305.14 0.32 305.645 ;
		RECT	0 306.935 0.32 307.72 ;
		RECT	0 308.02 0.32 308.525 ;
		RECT	0 309.815 0.32 310.6 ;
		RECT	0 310.9 0.32 311.405 ;
		RECT	0 312.695 0.32 313.48 ;
		RECT	0 313.78 0.32 314.285 ;
		RECT	0 315.575 0.32 316.36 ;
		RECT	0 316.66 0.32 317.165 ;
		RECT	0 318.455 0.32 319.24 ;
		RECT	0 319.54 0.32 320.045 ;
		RECT	0 321.335 0.32 322.12 ;
		RECT	0 322.42 0.32 322.925 ;
		RECT	0 324.215 0.32 325 ;
		RECT	0 325.3 0.32 325.805 ;
		RECT	0 327.095 0.32 327.88 ;
		RECT	0 328.18 0.32 328.685 ;
		RECT	0 329.975 0.32 330.76 ;
		RECT	0 331.06 0.32 331.565 ;
		RECT	0 332.855 0.32 333.64 ;
		RECT	0 333.94 0.32 334.445 ;
		RECT	0 335.735 0.32 336.52 ;
		RECT	0 336.82 0.32 337.325 ;
		RECT	0 338.615 0.32 339.4 ;
		RECT	0 339.7 0.32 340.205 ;
		RECT	0 341.495 0.32 342.28 ;
		RECT	0 342.58 0.32 343.085 ;
		RECT	0 344.375 0.32 345.16 ;
		RECT	0 345.46 0.32 345.965 ;
		RECT	0 347.255 0.32 348.04 ;
		RECT	0 348.34 0.32 348.845 ;
		RECT	0 350.135 0.32 350.92 ;
		RECT	0 351.22 0.32 351.725 ;
		RECT	0 353.015 0.32 353.8 ;
		RECT	0 354.1 0.32 354.605 ;
		RECT	0 355.895 0.32 356.68 ;
		RECT	0 356.98 0.32 357.485 ;
		RECT	0 358.775 0.32 359.56 ;
		RECT	0 359.86 0.32 360.365 ;
		RECT	0 361.655 0.32 362.44 ;
		RECT	0 362.74 0.32 363.245 ;
		RECT	0 364.535 0.32 365.32 ;
		RECT	0 365.62 0.32 366.125 ;
		RECT	0 367.415 0.32 368.2 ;
		RECT	0 368.5 0.32 369.005 ;
		RECT	0 370.295 0.32 371.08 ;
		RECT	0 371.38 0.32 371.885 ;
		RECT	0 373.175 0.32 373.96 ;
		RECT	0 374.26 0.32 374.765 ;
		RECT	0 376.055 0.32 376.84 ;
		RECT	0 377.14 0.32 377.645 ;
		RECT	0 378.935 0.32 379.72 ;
		RECT	0 380.02 0.32 380.525 ;
		RECT	0 381.815 0.32 382.6 ;
		RECT	0 382.9 0.32 383.405 ;
		RECT	0 384.695 0.32 385.48 ;
		RECT	0 385.78 0.32 386.285 ;
		RECT	0 387.575 0.32 388.36 ;
		RECT	0 388.66 0.32 389.165 ;
		RECT	0 390.455 0.32 391.24 ;
		RECT	0 391.54 0.32 392.045 ;
		RECT	0 393.335 0.32 394.12 ;
		RECT	0 394.42 0.32 394.925 ;
		RECT	0 396.215 0.32 397 ;
		RECT	0 397.3 0.32 397.805 ;
		RECT	0 399.095 0.32 399.88 ;
		RECT	0 400.18 0.32 400.685 ;
		RECT	0 401.975 0.32 402.76 ;
		RECT	0 403.06 0.32 403.565 ;
		RECT	0 404.855 0.32 405.64 ;
		RECT	0 405.94 0.32 406.445 ;
		RECT	0 407.735 0.32 408.52 ;
		RECT	0 408.82 0.32 409.325 ;
		RECT	0 410.615 0.32 411.4 ;
		RECT	0 411.7 0.32 412.205 ;
		RECT	0 413.495 0.32 414.3 ;
		RECT	21.655 0 21.975 414.86 ;
		RECT	0.32 0 21.655 0.35 ;
		RECT	0.32 414.51 21.655 414.86 ;
		LAYER	M2 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0.35 21.655 414.51 ;
		RECT	0 0.56 0.32 1.365 ;
		RECT	0 2.655 0.32 3.16 ;
		RECT	0 3.46 0.32 4.245 ;
		RECT	0 5.535 0.32 6.04 ;
		RECT	0 6.34 0.32 7.125 ;
		RECT	0 8.415 0.32 8.92 ;
		RECT	0 9.22 0.32 10.005 ;
		RECT	0 11.295 0.32 11.8 ;
		RECT	0 12.1 0.32 12.885 ;
		RECT	0 14.175 0.32 14.68 ;
		RECT	0 14.98 0.32 15.765 ;
		RECT	0 17.055 0.32 17.56 ;
		RECT	0 17.86 0.32 18.645 ;
		RECT	0 19.935 0.32 20.44 ;
		RECT	0 20.74 0.32 21.525 ;
		RECT	0 22.815 0.32 23.32 ;
		RECT	0 23.62 0.32 24.405 ;
		RECT	0 25.695 0.32 26.2 ;
		RECT	0 26.5 0.32 27.285 ;
		RECT	0 28.575 0.32 29.08 ;
		RECT	0 29.38 0.32 30.165 ;
		RECT	0 31.455 0.32 31.96 ;
		RECT	0 32.26 0.32 33.045 ;
		RECT	0 34.335 0.32 34.84 ;
		RECT	0 35.14 0.32 35.925 ;
		RECT	0 37.215 0.32 37.72 ;
		RECT	0 38.02 0.32 38.805 ;
		RECT	0 40.095 0.32 40.6 ;
		RECT	0 40.9 0.32 41.685 ;
		RECT	0 42.975 0.32 43.48 ;
		RECT	0 43.78 0.32 44.565 ;
		RECT	0 45.855 0.32 46.36 ;
		RECT	0 46.66 0.32 47.445 ;
		RECT	0 48.735 0.32 49.24 ;
		RECT	0 49.54 0.32 50.325 ;
		RECT	0 51.615 0.32 52.12 ;
		RECT	0 52.42 0.32 53.205 ;
		RECT	0 54.495 0.32 55 ;
		RECT	0 55.3 0.32 56.085 ;
		RECT	0 57.375 0.32 57.88 ;
		RECT	0 58.18 0.32 58.965 ;
		RECT	0 60.255 0.32 60.76 ;
		RECT	0 61.06 0.32 61.845 ;
		RECT	0 63.135 0.32 63.64 ;
		RECT	0 63.94 0.32 64.725 ;
		RECT	0 66.015 0.32 66.52 ;
		RECT	0 66.82 0.32 67.605 ;
		RECT	0 68.895 0.32 69.4 ;
		RECT	0 69.7 0.32 70.485 ;
		RECT	0 71.775 0.32 72.28 ;
		RECT	0 72.58 0.32 73.365 ;
		RECT	0 74.655 0.32 75.16 ;
		RECT	0 75.46 0.32 76.245 ;
		RECT	0 77.535 0.32 78.04 ;
		RECT	0 78.34 0.32 79.125 ;
		RECT	0 80.415 0.32 80.92 ;
		RECT	0 81.22 0.32 82.005 ;
		RECT	0 83.295 0.32 83.8 ;
		RECT	0 84.1 0.32 84.885 ;
		RECT	0 86.175 0.32 86.68 ;
		RECT	0 86.98 0.32 87.765 ;
		RECT	0 89.055 0.32 89.56 ;
		RECT	0 89.86 0.32 90.645 ;
		RECT	0 91.935 0.32 92.44 ;
		RECT	0 92.74 0.32 93.525 ;
		RECT	0 94.815 0.32 95.32 ;
		RECT	0 95.62 0.32 96.405 ;
		RECT	0 97.695 0.32 98.2 ;
		RECT	0 98.5 0.32 99.285 ;
		RECT	0 100.575 0.32 101.08 ;
		RECT	0 101.38 0.32 102.165 ;
		RECT	0 103.455 0.32 103.96 ;
		RECT	0 104.26 0.32 105.045 ;
		RECT	0 106.335 0.32 106.84 ;
		RECT	0 107.14 0.32 107.925 ;
		RECT	0 109.215 0.32 109.72 ;
		RECT	0 110.02 0.32 110.805 ;
		RECT	0 112.095 0.32 112.6 ;
		RECT	0 112.9 0.32 113.685 ;
		RECT	0 114.975 0.32 115.48 ;
		RECT	0 115.78 0.32 116.565 ;
		RECT	0 117.855 0.32 118.36 ;
		RECT	0 118.66 0.32 119.445 ;
		RECT	0 120.735 0.32 121.24 ;
		RECT	0 121.54 0.32 122.325 ;
		RECT	0 123.615 0.32 124.12 ;
		RECT	0 124.42 0.32 125.205 ;
		RECT	0 126.495 0.32 127 ;
		RECT	0 127.3 0.32 128.085 ;
		RECT	0 129.375 0.32 129.88 ;
		RECT	0 130.18 0.32 130.965 ;
		RECT	0 132.255 0.32 132.76 ;
		RECT	0 133.06 0.32 133.845 ;
		RECT	0 135.135 0.32 135.64 ;
		RECT	0 135.94 0.32 136.725 ;
		RECT	0 138.015 0.32 138.52 ;
		RECT	0 138.82 0.32 139.605 ;
		RECT	0 140.895 0.32 141.4 ;
		RECT	0 141.7 0.32 142.485 ;
		RECT	0 143.775 0.32 144.28 ;
		RECT	0 144.58 0.32 145.365 ;
		RECT	0 146.655 0.32 147.16 ;
		RECT	0 147.46 0.32 148.245 ;
		RECT	0 149.535 0.32 150.04 ;
		RECT	0 150.34 0.32 151.125 ;
		RECT	0 152.415 0.32 152.92 ;
		RECT	0 153.22 0.32 154.005 ;
		RECT	0 155.295 0.32 155.8 ;
		RECT	0 156.1 0.32 156.885 ;
		RECT	0 158.175 0.32 158.68 ;
		RECT	0 158.98 0.32 159.765 ;
		RECT	0 161.055 0.32 161.56 ;
		RECT	0 161.86 0.32 162.645 ;
		RECT	0 163.935 0.32 164.44 ;
		RECT	0 164.74 0.32 165.525 ;
		RECT	0 166.815 0.32 167.32 ;
		RECT	0 167.62 0.32 168.405 ;
		RECT	0 169.695 0.32 170.2 ;
		RECT	0 170.5 0.32 171.285 ;
		RECT	0 172.575 0.32 173.08 ;
		RECT	0 173.38 0.32 174.165 ;
		RECT	0 175.455 0.32 175.96 ;
		RECT	0 176.26 0.32 177.045 ;
		RECT	0 178.335 0.32 178.84 ;
		RECT	0 179.14 0.32 179.925 ;
		RECT	0 181.215 0.32 181.72 ;
		RECT	0 182.02 0.32 182.805 ;
		RECT	0 184.095 0.32 184.6 ;
		RECT	0 184.9 0.32 187 ;
		RECT	0 187.3 0.32 187.35 ;
		RECT	0 187.65 0.32 188.01 ;
		RECT	0 188.71 0.32 190.35 ;
		RECT	0 190.955 0.32 191.17 ;
		RECT	0 191.47 0.32 191.575 ;
		RECT	0 191.875 0.32 193.685 ;
		RECT	0 193.985 0.32 194.2 ;
		RECT	0 194.5 0.32 194.605 ;
		RECT	0 194.905 0.32 196.745 ;
		RECT	0 197.045 0.32 197.23 ;
		RECT	0 197.53 0.32 197.635 ;
		RECT	0 197.935 0.32 198.03 ;
		RECT	0 198.33 0.32 198.4 ;
		RECT	0 198.7 0.32 198.775 ;
		RECT	0 199.075 0.32 199.26 ;
		RECT	0 199.97 0.32 201.405 ;
		RECT	0 202.105 0.32 202.29 ;
		RECT	0 202.875 0.32 205.8 ;
		RECT	0 206.5 0.32 206.97 ;
		RECT	0 207.27 0.32 208.635 ;
		RECT	0 208.935 0.32 212.725 ;
		RECT	0 213.26 0.32 213.45 ;
		RECT	0 213.75 0.32 213.825 ;
		RECT	0 214.125 0.32 214.205 ;
		RECT	0 214.505 0.32 215.205 ;
		RECT	0 215.505 0.32 215.995 ;
		RECT	0 216.295 0.32 216.48 ;
		RECT	0 216.78 0.32 216.885 ;
		RECT	0 217.185 0.32 217.65 ;
		RECT	0 217.95 0.32 218.025 ;
		RECT	0 218.325 0.32 218.48 ;
		RECT	0 218.98 0.32 220.225 ;
		RECT	0 220.525 0.32 220.65 ;
		RECT	0 221.16 0.32 221.54 ;
		RECT	0 221.84 0.32 223.68 ;
		RECT	0 223.98 0.32 224.085 ;
		RECT	0 224.385 0.32 224.57 ;
		RECT	0 225.125 0.32 225.6 ;
		RECT	0 225.9 0.32 228.21 ;
		RECT	0 228.51 0.32 228.605 ;
		RECT	0 228.905 0.32 229.15 ;
		RECT	0 229.45 0.32 229.96 ;
		RECT	0 230.26 0.32 230.765 ;
		RECT	0 232.055 0.32 232.84 ;
		RECT	0 233.14 0.32 233.645 ;
		RECT	0 234.935 0.32 235.72 ;
		RECT	0 236.02 0.32 236.525 ;
		RECT	0 237.815 0.32 238.6 ;
		RECT	0 238.9 0.32 239.405 ;
		RECT	0 240.695 0.32 241.48 ;
		RECT	0 241.78 0.32 242.285 ;
		RECT	0 243.575 0.32 244.36 ;
		RECT	0 244.66 0.32 245.165 ;
		RECT	0 246.455 0.32 247.24 ;
		RECT	0 247.54 0.32 248.045 ;
		RECT	0 249.335 0.32 250.12 ;
		RECT	0 250.42 0.32 250.925 ;
		RECT	0 252.215 0.32 253 ;
		RECT	0 253.3 0.32 253.805 ;
		RECT	0 255.095 0.32 255.88 ;
		RECT	0 256.18 0.32 256.685 ;
		RECT	0 257.975 0.32 258.76 ;
		RECT	0 259.06 0.32 259.565 ;
		RECT	0 260.855 0.32 261.64 ;
		RECT	0 261.94 0.32 262.445 ;
		RECT	0 263.735 0.32 264.52 ;
		RECT	0 264.82 0.32 265.325 ;
		RECT	0 266.615 0.32 267.4 ;
		RECT	0 267.7 0.32 268.205 ;
		RECT	0 269.495 0.32 270.28 ;
		RECT	0 270.58 0.32 271.085 ;
		RECT	0 272.375 0.32 273.16 ;
		RECT	0 273.46 0.32 273.965 ;
		RECT	0 275.255 0.32 276.04 ;
		RECT	0 276.34 0.32 276.845 ;
		RECT	0 278.135 0.32 278.92 ;
		RECT	0 279.22 0.32 279.725 ;
		RECT	0 281.015 0.32 281.8 ;
		RECT	0 282.1 0.32 282.605 ;
		RECT	0 283.895 0.32 284.68 ;
		RECT	0 284.98 0.32 285.485 ;
		RECT	0 286.775 0.32 287.56 ;
		RECT	0 287.86 0.32 288.365 ;
		RECT	0 289.655 0.32 290.44 ;
		RECT	0 290.74 0.32 291.245 ;
		RECT	0 292.535 0.32 293.32 ;
		RECT	0 293.62 0.32 294.125 ;
		RECT	0 295.415 0.32 296.2 ;
		RECT	0 296.5 0.32 297.005 ;
		RECT	0 298.295 0.32 299.08 ;
		RECT	0 299.38 0.32 299.885 ;
		RECT	0 301.175 0.32 301.96 ;
		RECT	0 302.26 0.32 302.765 ;
		RECT	0 304.055 0.32 304.84 ;
		RECT	0 305.14 0.32 305.645 ;
		RECT	0 306.935 0.32 307.72 ;
		RECT	0 308.02 0.32 308.525 ;
		RECT	0 309.815 0.32 310.6 ;
		RECT	0 310.9 0.32 311.405 ;
		RECT	0 312.695 0.32 313.48 ;
		RECT	0 313.78 0.32 314.285 ;
		RECT	0 315.575 0.32 316.36 ;
		RECT	0 316.66 0.32 317.165 ;
		RECT	0 318.455 0.32 319.24 ;
		RECT	0 319.54 0.32 320.045 ;
		RECT	0 321.335 0.32 322.12 ;
		RECT	0 322.42 0.32 322.925 ;
		RECT	0 324.215 0.32 325 ;
		RECT	0 325.3 0.32 325.805 ;
		RECT	0 327.095 0.32 327.88 ;
		RECT	0 328.18 0.32 328.685 ;
		RECT	0 329.975 0.32 330.76 ;
		RECT	0 331.06 0.32 331.565 ;
		RECT	0 332.855 0.32 333.64 ;
		RECT	0 333.94 0.32 334.445 ;
		RECT	0 335.735 0.32 336.52 ;
		RECT	0 336.82 0.32 337.325 ;
		RECT	0 338.615 0.32 339.4 ;
		RECT	0 339.7 0.32 340.205 ;
		RECT	0 341.495 0.32 342.28 ;
		RECT	0 342.58 0.32 343.085 ;
		RECT	0 344.375 0.32 345.16 ;
		RECT	0 345.46 0.32 345.965 ;
		RECT	0 347.255 0.32 348.04 ;
		RECT	0 348.34 0.32 348.845 ;
		RECT	0 350.135 0.32 350.92 ;
		RECT	0 351.22 0.32 351.725 ;
		RECT	0 353.015 0.32 353.8 ;
		RECT	0 354.1 0.32 354.605 ;
		RECT	0 355.895 0.32 356.68 ;
		RECT	0 356.98 0.32 357.485 ;
		RECT	0 358.775 0.32 359.56 ;
		RECT	0 359.86 0.32 360.365 ;
		RECT	0 361.655 0.32 362.44 ;
		RECT	0 362.74 0.32 363.245 ;
		RECT	0 364.535 0.32 365.32 ;
		RECT	0 365.62 0.32 366.125 ;
		RECT	0 367.415 0.32 368.2 ;
		RECT	0 368.5 0.32 369.005 ;
		RECT	0 370.295 0.32 371.08 ;
		RECT	0 371.38 0.32 371.885 ;
		RECT	0 373.175 0.32 373.96 ;
		RECT	0 374.26 0.32 374.765 ;
		RECT	0 376.055 0.32 376.84 ;
		RECT	0 377.14 0.32 377.645 ;
		RECT	0 378.935 0.32 379.72 ;
		RECT	0 380.02 0.32 380.525 ;
		RECT	0 381.815 0.32 382.6 ;
		RECT	0 382.9 0.32 383.405 ;
		RECT	0 384.695 0.32 385.48 ;
		RECT	0 385.78 0.32 386.285 ;
		RECT	0 387.575 0.32 388.36 ;
		RECT	0 388.66 0.32 389.165 ;
		RECT	0 390.455 0.32 391.24 ;
		RECT	0 391.54 0.32 392.045 ;
		RECT	0 393.335 0.32 394.12 ;
		RECT	0 394.42 0.32 394.925 ;
		RECT	0 396.215 0.32 397 ;
		RECT	0 397.3 0.32 397.805 ;
		RECT	0 399.095 0.32 399.88 ;
		RECT	0 400.18 0.32 400.685 ;
		RECT	0 401.975 0.32 402.76 ;
		RECT	0 403.06 0.32 403.565 ;
		RECT	0 404.855 0.32 405.64 ;
		RECT	0 405.94 0.32 406.445 ;
		RECT	0 407.735 0.32 408.52 ;
		RECT	0 408.82 0.32 409.325 ;
		RECT	0 410.615 0.32 411.4 ;
		RECT	0 411.7 0.32 412.205 ;
		RECT	0 413.495 0.32 414.3 ;
		RECT	21.655 0 21.975 414.86 ;
		RECT	0.32 0 21.655 0.35 ;
		RECT	0.32 414.51 21.655 414.86 ;
		LAYER	M3 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0.35 21.655 414.51 ;
		RECT	0 0.56 0.32 1.365 ;
		RECT	0 2.655 0.32 3.16 ;
		RECT	0 3.46 0.32 4.245 ;
		RECT	0 5.535 0.32 6.04 ;
		RECT	0 6.34 0.32 7.125 ;
		RECT	0 8.415 0.32 8.92 ;
		RECT	0 9.22 0.32 10.005 ;
		RECT	0 11.295 0.32 11.8 ;
		RECT	0 12.1 0.32 12.885 ;
		RECT	0 14.175 0.32 14.68 ;
		RECT	0 14.98 0.32 15.765 ;
		RECT	0 17.055 0.32 17.56 ;
		RECT	0 17.86 0.32 18.645 ;
		RECT	0 19.935 0.32 20.44 ;
		RECT	0 20.74 0.32 21.525 ;
		RECT	0 22.815 0.32 23.32 ;
		RECT	0 23.62 0.32 24.405 ;
		RECT	0 25.695 0.32 26.2 ;
		RECT	0 26.5 0.32 27.285 ;
		RECT	0 28.575 0.32 29.08 ;
		RECT	0 29.38 0.32 30.165 ;
		RECT	0 31.455 0.32 31.96 ;
		RECT	0 32.26 0.32 33.045 ;
		RECT	0 34.335 0.32 34.84 ;
		RECT	0 35.14 0.32 35.925 ;
		RECT	0 37.215 0.32 37.72 ;
		RECT	0 38.02 0.32 38.805 ;
		RECT	0 40.095 0.32 40.6 ;
		RECT	0 40.9 0.32 41.685 ;
		RECT	0 42.975 0.32 43.48 ;
		RECT	0 43.78 0.32 44.565 ;
		RECT	0 45.855 0.32 46.36 ;
		RECT	0 46.66 0.32 47.445 ;
		RECT	0 48.735 0.32 49.24 ;
		RECT	0 49.54 0.32 50.325 ;
		RECT	0 51.615 0.32 52.12 ;
		RECT	0 52.42 0.32 53.205 ;
		RECT	0 54.495 0.32 55 ;
		RECT	0 55.3 0.32 56.085 ;
		RECT	0 57.375 0.32 57.88 ;
		RECT	0 58.18 0.32 58.965 ;
		RECT	0 60.255 0.32 60.76 ;
		RECT	0 61.06 0.32 61.845 ;
		RECT	0 63.135 0.32 63.64 ;
		RECT	0 63.94 0.32 64.725 ;
		RECT	0 66.015 0.32 66.52 ;
		RECT	0 66.82 0.32 67.605 ;
		RECT	0 68.895 0.32 69.4 ;
		RECT	0 69.7 0.32 70.485 ;
		RECT	0 71.775 0.32 72.28 ;
		RECT	0 72.58 0.32 73.365 ;
		RECT	0 74.655 0.32 75.16 ;
		RECT	0 75.46 0.32 76.245 ;
		RECT	0 77.535 0.32 78.04 ;
		RECT	0 78.34 0.32 79.125 ;
		RECT	0 80.415 0.32 80.92 ;
		RECT	0 81.22 0.32 82.005 ;
		RECT	0 83.295 0.32 83.8 ;
		RECT	0 84.1 0.32 84.885 ;
		RECT	0 86.175 0.32 86.68 ;
		RECT	0 86.98 0.32 87.765 ;
		RECT	0 89.055 0.32 89.56 ;
		RECT	0 89.86 0.32 90.645 ;
		RECT	0 91.935 0.32 92.44 ;
		RECT	0 92.74 0.32 93.525 ;
		RECT	0 94.815 0.32 95.32 ;
		RECT	0 95.62 0.32 96.405 ;
		RECT	0 97.695 0.32 98.2 ;
		RECT	0 98.5 0.32 99.285 ;
		RECT	0 100.575 0.32 101.08 ;
		RECT	0 101.38 0.32 102.165 ;
		RECT	0 103.455 0.32 103.96 ;
		RECT	0 104.26 0.32 105.045 ;
		RECT	0 106.335 0.32 106.84 ;
		RECT	0 107.14 0.32 107.925 ;
		RECT	0 109.215 0.32 109.72 ;
		RECT	0 110.02 0.32 110.805 ;
		RECT	0 112.095 0.32 112.6 ;
		RECT	0 112.9 0.32 113.685 ;
		RECT	0 114.975 0.32 115.48 ;
		RECT	0 115.78 0.32 116.565 ;
		RECT	0 117.855 0.32 118.36 ;
		RECT	0 118.66 0.32 119.445 ;
		RECT	0 120.735 0.32 121.24 ;
		RECT	0 121.54 0.32 122.325 ;
		RECT	0 123.615 0.32 124.12 ;
		RECT	0 124.42 0.32 125.205 ;
		RECT	0 126.495 0.32 127 ;
		RECT	0 127.3 0.32 128.085 ;
		RECT	0 129.375 0.32 129.88 ;
		RECT	0 130.18 0.32 130.965 ;
		RECT	0 132.255 0.32 132.76 ;
		RECT	0 133.06 0.32 133.845 ;
		RECT	0 135.135 0.32 135.64 ;
		RECT	0 135.94 0.32 136.725 ;
		RECT	0 138.015 0.32 138.52 ;
		RECT	0 138.82 0.32 139.605 ;
		RECT	0 140.895 0.32 141.4 ;
		RECT	0 141.7 0.32 142.485 ;
		RECT	0 143.775 0.32 144.28 ;
		RECT	0 144.58 0.32 145.365 ;
		RECT	0 146.655 0.32 147.16 ;
		RECT	0 147.46 0.32 148.245 ;
		RECT	0 149.535 0.32 150.04 ;
		RECT	0 150.34 0.32 151.125 ;
		RECT	0 152.415 0.32 152.92 ;
		RECT	0 153.22 0.32 154.005 ;
		RECT	0 155.295 0.32 155.8 ;
		RECT	0 156.1 0.32 156.885 ;
		RECT	0 158.175 0.32 158.68 ;
		RECT	0 158.98 0.32 159.765 ;
		RECT	0 161.055 0.32 161.56 ;
		RECT	0 161.86 0.32 162.645 ;
		RECT	0 163.935 0.32 164.44 ;
		RECT	0 164.74 0.32 165.525 ;
		RECT	0 166.815 0.32 167.32 ;
		RECT	0 167.62 0.32 168.405 ;
		RECT	0 169.695 0.32 170.2 ;
		RECT	0 170.5 0.32 171.285 ;
		RECT	0 172.575 0.32 173.08 ;
		RECT	0 173.38 0.32 174.165 ;
		RECT	0 175.455 0.32 175.96 ;
		RECT	0 176.26 0.32 177.045 ;
		RECT	0 178.335 0.32 178.84 ;
		RECT	0 179.14 0.32 179.925 ;
		RECT	0 181.215 0.32 181.72 ;
		RECT	0 182.02 0.32 182.805 ;
		RECT	0 184.095 0.32 184.6 ;
		RECT	0 184.9 0.32 187 ;
		RECT	0 187.3 0.32 187.35 ;
		RECT	0 187.65 0.32 188.01 ;
		RECT	0 188.71 0.32 190.35 ;
		RECT	0 190.955 0.32 191.17 ;
		RECT	0 191.47 0.32 191.575 ;
		RECT	0 191.875 0.32 193.685 ;
		RECT	0 193.985 0.32 194.2 ;
		RECT	0 194.5 0.32 194.605 ;
		RECT	0 194.905 0.32 196.745 ;
		RECT	0 197.045 0.32 197.23 ;
		RECT	0 197.53 0.32 197.635 ;
		RECT	0 197.935 0.32 198.03 ;
		RECT	0 198.33 0.32 198.4 ;
		RECT	0 198.7 0.32 198.775 ;
		RECT	0 199.075 0.32 199.26 ;
		RECT	0 199.97 0.32 201.405 ;
		RECT	0 202.105 0.32 202.29 ;
		RECT	0 202.875 0.32 205.8 ;
		RECT	0 206.5 0.32 206.97 ;
		RECT	0 207.27 0.32 208.635 ;
		RECT	0 208.935 0.32 212.725 ;
		RECT	0 213.26 0.32 213.45 ;
		RECT	0 213.75 0.32 213.825 ;
		RECT	0 214.125 0.32 214.205 ;
		RECT	0 214.505 0.32 215.205 ;
		RECT	0 215.505 0.32 215.995 ;
		RECT	0 216.295 0.32 216.48 ;
		RECT	0 216.78 0.32 216.885 ;
		RECT	0 217.185 0.32 217.65 ;
		RECT	0 217.95 0.32 218.025 ;
		RECT	0 218.325 0.32 218.48 ;
		RECT	0 218.98 0.32 220.225 ;
		RECT	0 220.525 0.32 220.65 ;
		RECT	0 221.16 0.32 221.54 ;
		RECT	0 221.84 0.32 223.68 ;
		RECT	0 223.98 0.32 224.085 ;
		RECT	0 224.385 0.32 224.57 ;
		RECT	0 225.125 0.32 225.6 ;
		RECT	0 225.9 0.32 228.21 ;
		RECT	0 228.51 0.32 228.605 ;
		RECT	0 228.905 0.32 229.15 ;
		RECT	0 229.45 0.32 229.96 ;
		RECT	0 230.26 0.32 230.765 ;
		RECT	0 232.055 0.32 232.84 ;
		RECT	0 233.14 0.32 233.645 ;
		RECT	0 234.935 0.32 235.72 ;
		RECT	0 236.02 0.32 236.525 ;
		RECT	0 237.815 0.32 238.6 ;
		RECT	0 238.9 0.32 239.405 ;
		RECT	0 240.695 0.32 241.48 ;
		RECT	0 241.78 0.32 242.285 ;
		RECT	0 243.575 0.32 244.36 ;
		RECT	0 244.66 0.32 245.165 ;
		RECT	0 246.455 0.32 247.24 ;
		RECT	0 247.54 0.32 248.045 ;
		RECT	0 249.335 0.32 250.12 ;
		RECT	0 250.42 0.32 250.925 ;
		RECT	0 252.215 0.32 253 ;
		RECT	0 253.3 0.32 253.805 ;
		RECT	0 255.095 0.32 255.88 ;
		RECT	0 256.18 0.32 256.685 ;
		RECT	0 257.975 0.32 258.76 ;
		RECT	0 259.06 0.32 259.565 ;
		RECT	0 260.855 0.32 261.64 ;
		RECT	0 261.94 0.32 262.445 ;
		RECT	0 263.735 0.32 264.52 ;
		RECT	0 264.82 0.32 265.325 ;
		RECT	0 266.615 0.32 267.4 ;
		RECT	0 267.7 0.32 268.205 ;
		RECT	0 269.495 0.32 270.28 ;
		RECT	0 270.58 0.32 271.085 ;
		RECT	0 272.375 0.32 273.16 ;
		RECT	0 273.46 0.32 273.965 ;
		RECT	0 275.255 0.32 276.04 ;
		RECT	0 276.34 0.32 276.845 ;
		RECT	0 278.135 0.32 278.92 ;
		RECT	0 279.22 0.32 279.725 ;
		RECT	0 281.015 0.32 281.8 ;
		RECT	0 282.1 0.32 282.605 ;
		RECT	0 283.895 0.32 284.68 ;
		RECT	0 284.98 0.32 285.485 ;
		RECT	0 286.775 0.32 287.56 ;
		RECT	0 287.86 0.32 288.365 ;
		RECT	0 289.655 0.32 290.44 ;
		RECT	0 290.74 0.32 291.245 ;
		RECT	0 292.535 0.32 293.32 ;
		RECT	0 293.62 0.32 294.125 ;
		RECT	0 295.415 0.32 296.2 ;
		RECT	0 296.5 0.32 297.005 ;
		RECT	0 298.295 0.32 299.08 ;
		RECT	0 299.38 0.32 299.885 ;
		RECT	0 301.175 0.32 301.96 ;
		RECT	0 302.26 0.32 302.765 ;
		RECT	0 304.055 0.32 304.84 ;
		RECT	0 305.14 0.32 305.645 ;
		RECT	0 306.935 0.32 307.72 ;
		RECT	0 308.02 0.32 308.525 ;
		RECT	0 309.815 0.32 310.6 ;
		RECT	0 310.9 0.32 311.405 ;
		RECT	0 312.695 0.32 313.48 ;
		RECT	0 313.78 0.32 314.285 ;
		RECT	0 315.575 0.32 316.36 ;
		RECT	0 316.66 0.32 317.165 ;
		RECT	0 318.455 0.32 319.24 ;
		RECT	0 319.54 0.32 320.045 ;
		RECT	0 321.335 0.32 322.12 ;
		RECT	0 322.42 0.32 322.925 ;
		RECT	0 324.215 0.32 325 ;
		RECT	0 325.3 0.32 325.805 ;
		RECT	0 327.095 0.32 327.88 ;
		RECT	0 328.18 0.32 328.685 ;
		RECT	0 329.975 0.32 330.76 ;
		RECT	0 331.06 0.32 331.565 ;
		RECT	0 332.855 0.32 333.64 ;
		RECT	0 333.94 0.32 334.445 ;
		RECT	0 335.735 0.32 336.52 ;
		RECT	0 336.82 0.32 337.325 ;
		RECT	0 338.615 0.32 339.4 ;
		RECT	0 339.7 0.32 340.205 ;
		RECT	0 341.495 0.32 342.28 ;
		RECT	0 342.58 0.32 343.085 ;
		RECT	0 344.375 0.32 345.16 ;
		RECT	0 345.46 0.32 345.965 ;
		RECT	0 347.255 0.32 348.04 ;
		RECT	0 348.34 0.32 348.845 ;
		RECT	0 350.135 0.32 350.92 ;
		RECT	0 351.22 0.32 351.725 ;
		RECT	0 353.015 0.32 353.8 ;
		RECT	0 354.1 0.32 354.605 ;
		RECT	0 355.895 0.32 356.68 ;
		RECT	0 356.98 0.32 357.485 ;
		RECT	0 358.775 0.32 359.56 ;
		RECT	0 359.86 0.32 360.365 ;
		RECT	0 361.655 0.32 362.44 ;
		RECT	0 362.74 0.32 363.245 ;
		RECT	0 364.535 0.32 365.32 ;
		RECT	0 365.62 0.32 366.125 ;
		RECT	0 367.415 0.32 368.2 ;
		RECT	0 368.5 0.32 369.005 ;
		RECT	0 370.295 0.32 371.08 ;
		RECT	0 371.38 0.32 371.885 ;
		RECT	0 373.175 0.32 373.96 ;
		RECT	0 374.26 0.32 374.765 ;
		RECT	0 376.055 0.32 376.84 ;
		RECT	0 377.14 0.32 377.645 ;
		RECT	0 378.935 0.32 379.72 ;
		RECT	0 380.02 0.32 380.525 ;
		RECT	0 381.815 0.32 382.6 ;
		RECT	0 382.9 0.32 383.405 ;
		RECT	0 384.695 0.32 385.48 ;
		RECT	0 385.78 0.32 386.285 ;
		RECT	0 387.575 0.32 388.36 ;
		RECT	0 388.66 0.32 389.165 ;
		RECT	0 390.455 0.32 391.24 ;
		RECT	0 391.54 0.32 392.045 ;
		RECT	0 393.335 0.32 394.12 ;
		RECT	0 394.42 0.32 394.925 ;
		RECT	0 396.215 0.32 397 ;
		RECT	0 397.3 0.32 397.805 ;
		RECT	0 399.095 0.32 399.88 ;
		RECT	0 400.18 0.32 400.685 ;
		RECT	0 401.975 0.32 402.76 ;
		RECT	0 403.06 0.32 403.565 ;
		RECT	0 404.855 0.32 405.64 ;
		RECT	0 405.94 0.32 406.445 ;
		RECT	0 407.735 0.32 408.52 ;
		RECT	0 408.82 0.32 409.325 ;
		RECT	0 410.615 0.32 411.4 ;
		RECT	0 411.7 0.32 412.205 ;
		RECT	0 413.495 0.32 414.3 ;
		RECT	21.655 0 21.975 414.86 ;
		RECT	0.32 0 21.655 0.35 ;
		RECT	0.32 414.51 21.655 414.86 ;
		LAYER	M4 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0 21.655 0.105 ;
		RECT	0 0 0.32 0.105 ;
		RECT	21.655 0 21.975 0.105 ;
		RECT	0.32 1.335 21.655 1.885 ;
		RECT	0 1.335 0.32 1.885 ;
		RECT	21.655 1.335 21.975 1.885 ;
		RECT	0.32 2.435 21.655 3.215 ;
		RECT	0 2.435 0.32 3.215 ;
		RECT	21.655 2.435 21.975 3.215 ;
		RECT	0.32 4.215 21.655 4.765 ;
		RECT	0 4.215 0.32 4.765 ;
		RECT	21.655 4.215 21.975 4.765 ;
		RECT	0.32 5.315 21.655 6.095 ;
		RECT	0 5.315 0.32 6.095 ;
		RECT	21.655 5.315 21.975 6.095 ;
		RECT	0.32 7.095 21.655 7.645 ;
		RECT	0 7.095 0.32 7.645 ;
		RECT	21.655 7.095 21.975 7.645 ;
		RECT	0.32 8.195 21.655 8.975 ;
		RECT	0 8.195 0.32 8.975 ;
		RECT	21.655 8.195 21.975 8.975 ;
		RECT	0.32 9.975 21.655 10.525 ;
		RECT	0 9.975 0.32 10.525 ;
		RECT	21.655 9.975 21.975 10.525 ;
		RECT	0.32 11.075 21.655 11.855 ;
		RECT	0 11.075 0.32 11.855 ;
		RECT	21.655 11.075 21.975 11.855 ;
		RECT	0.32 12.855 21.655 13.405 ;
		RECT	0 12.855 0.32 13.405 ;
		RECT	21.655 12.855 21.975 13.405 ;
		RECT	0.32 13.955 21.655 14.735 ;
		RECT	0 13.955 0.32 14.735 ;
		RECT	21.655 13.955 21.975 14.735 ;
		RECT	0.32 15.735 21.655 16.285 ;
		RECT	0 15.735 0.32 16.285 ;
		RECT	21.655 15.735 21.975 16.285 ;
		RECT	0.32 16.835 21.655 17.615 ;
		RECT	0 16.835 0.32 17.615 ;
		RECT	21.655 16.835 21.975 17.615 ;
		RECT	0.32 18.615 21.655 19.165 ;
		RECT	0 18.615 0.32 19.165 ;
		RECT	21.655 18.615 21.975 19.165 ;
		RECT	0.32 19.715 21.655 20.495 ;
		RECT	0 19.715 0.32 20.495 ;
		RECT	21.655 19.715 21.975 20.495 ;
		RECT	0.32 21.495 21.655 22.045 ;
		RECT	0 21.495 0.32 22.045 ;
		RECT	21.655 21.495 21.975 22.045 ;
		RECT	0.32 22.595 21.655 23.375 ;
		RECT	0 22.595 0.32 23.375 ;
		RECT	21.655 22.595 21.975 23.375 ;
		RECT	0.32 24.375 21.655 24.925 ;
		RECT	0 24.375 0.32 24.925 ;
		RECT	21.655 24.375 21.975 24.925 ;
		RECT	0.32 25.475 21.655 26.255 ;
		RECT	0 25.475 0.32 26.255 ;
		RECT	21.655 25.475 21.975 26.255 ;
		RECT	0.32 27.255 21.655 27.805 ;
		RECT	0 27.255 0.32 27.805 ;
		RECT	21.655 27.255 21.975 27.805 ;
		RECT	0.32 28.355 21.655 29.135 ;
		RECT	0 28.355 0.32 29.135 ;
		RECT	21.655 28.355 21.975 29.135 ;
		RECT	0.32 30.135 21.655 30.685 ;
		RECT	0 30.135 0.32 30.685 ;
		RECT	21.655 30.135 21.975 30.685 ;
		RECT	0.32 31.235 21.655 32.015 ;
		RECT	0 31.235 0.32 32.015 ;
		RECT	21.655 31.235 21.975 32.015 ;
		RECT	0.32 33.015 21.655 33.565 ;
		RECT	0 33.015 0.32 33.565 ;
		RECT	21.655 33.015 21.975 33.565 ;
		RECT	0.32 34.115 21.655 34.895 ;
		RECT	0 34.115 0.32 34.895 ;
		RECT	21.655 34.115 21.975 34.895 ;
		RECT	0.32 35.895 21.655 36.445 ;
		RECT	0 35.895 0.32 36.445 ;
		RECT	21.655 35.895 21.975 36.445 ;
		RECT	0.32 36.995 21.655 37.775 ;
		RECT	0 36.995 0.32 37.775 ;
		RECT	21.655 36.995 21.975 37.775 ;
		RECT	0.32 38.775 21.655 39.325 ;
		RECT	0 38.775 0.32 39.325 ;
		RECT	21.655 38.775 21.975 39.325 ;
		RECT	0.32 39.875 21.655 40.655 ;
		RECT	0 39.875 0.32 40.655 ;
		RECT	21.655 39.875 21.975 40.655 ;
		RECT	0.32 41.655 21.655 42.205 ;
		RECT	0 41.655 0.32 42.205 ;
		RECT	21.655 41.655 21.975 42.205 ;
		RECT	0.32 42.755 21.655 43.535 ;
		RECT	0 42.755 0.32 43.535 ;
		RECT	21.655 42.755 21.975 43.535 ;
		RECT	0.32 44.535 21.655 45.085 ;
		RECT	0 44.535 0.32 45.085 ;
		RECT	21.655 44.535 21.975 45.085 ;
		RECT	0.32 45.635 21.655 46.415 ;
		RECT	0 45.635 0.32 46.415 ;
		RECT	21.655 45.635 21.975 46.415 ;
		RECT	0.32 47.415 21.655 47.965 ;
		RECT	0 47.415 0.32 47.965 ;
		RECT	21.655 47.415 21.975 47.965 ;
		RECT	0.32 48.515 21.655 49.295 ;
		RECT	0 48.515 0.32 49.295 ;
		RECT	21.655 48.515 21.975 49.295 ;
		RECT	0.32 50.295 21.655 50.845 ;
		RECT	0 50.295 0.32 50.845 ;
		RECT	21.655 50.295 21.975 50.845 ;
		RECT	0.32 51.395 21.655 52.175 ;
		RECT	0 51.395 0.32 52.175 ;
		RECT	21.655 51.395 21.975 52.175 ;
		RECT	0.32 53.175 21.655 53.725 ;
		RECT	0 53.175 0.32 53.725 ;
		RECT	21.655 53.175 21.975 53.725 ;
		RECT	0.32 54.275 21.655 55.055 ;
		RECT	0 54.275 0.32 55.055 ;
		RECT	21.655 54.275 21.975 55.055 ;
		RECT	0.32 56.055 21.655 56.605 ;
		RECT	0 56.055 0.32 56.605 ;
		RECT	21.655 56.055 21.975 56.605 ;
		RECT	0.32 57.155 21.655 57.935 ;
		RECT	0 57.155 0.32 57.935 ;
		RECT	21.655 57.155 21.975 57.935 ;
		RECT	0.32 58.935 21.655 59.485 ;
		RECT	0 58.935 0.32 59.485 ;
		RECT	21.655 58.935 21.975 59.485 ;
		RECT	0.32 60.035 21.655 60.815 ;
		RECT	0 60.035 0.32 60.815 ;
		RECT	21.655 60.035 21.975 60.815 ;
		RECT	0.32 61.815 21.655 62.365 ;
		RECT	0 61.815 0.32 62.365 ;
		RECT	21.655 61.815 21.975 62.365 ;
		RECT	0.32 62.915 21.655 63.695 ;
		RECT	0 62.915 0.32 63.695 ;
		RECT	21.655 62.915 21.975 63.695 ;
		RECT	0.32 64.695 21.655 65.245 ;
		RECT	0 64.695 0.32 65.245 ;
		RECT	21.655 64.695 21.975 65.245 ;
		RECT	0.32 65.795 21.655 66.575 ;
		RECT	0 65.795 0.32 66.575 ;
		RECT	21.655 65.795 21.975 66.575 ;
		RECT	0.32 67.575 21.655 68.125 ;
		RECT	0 67.575 0.32 68.125 ;
		RECT	21.655 67.575 21.975 68.125 ;
		RECT	0.32 68.675 21.655 69.455 ;
		RECT	0 68.675 0.32 69.455 ;
		RECT	21.655 68.675 21.975 69.455 ;
		RECT	0.32 70.455 21.655 71.005 ;
		RECT	0 70.455 0.32 71.005 ;
		RECT	21.655 70.455 21.975 71.005 ;
		RECT	0.32 71.555 21.655 72.335 ;
		RECT	0 71.555 0.32 72.335 ;
		RECT	21.655 71.555 21.975 72.335 ;
		RECT	0.32 73.335 21.655 73.885 ;
		RECT	0 73.335 0.32 73.885 ;
		RECT	21.655 73.335 21.975 73.885 ;
		RECT	0.32 74.435 21.655 75.215 ;
		RECT	0 74.435 0.32 75.215 ;
		RECT	21.655 74.435 21.975 75.215 ;
		RECT	0.32 76.215 21.655 76.765 ;
		RECT	0 76.215 0.32 76.765 ;
		RECT	21.655 76.215 21.975 76.765 ;
		RECT	0.32 77.315 21.655 78.095 ;
		RECT	0 77.315 0.32 78.095 ;
		RECT	21.655 77.315 21.975 78.095 ;
		RECT	0.32 79.095 21.655 79.645 ;
		RECT	0 79.095 0.32 79.645 ;
		RECT	21.655 79.095 21.975 79.645 ;
		RECT	0.32 80.195 21.655 80.975 ;
		RECT	0 80.195 0.32 80.975 ;
		RECT	21.655 80.195 21.975 80.975 ;
		RECT	0.32 81.975 21.655 82.525 ;
		RECT	0 81.975 0.32 82.525 ;
		RECT	21.655 81.975 21.975 82.525 ;
		RECT	0.32 83.075 21.655 83.855 ;
		RECT	0 83.075 0.32 83.855 ;
		RECT	21.655 83.075 21.975 83.855 ;
		RECT	0.32 84.855 21.655 85.405 ;
		RECT	0 84.855 0.32 85.405 ;
		RECT	21.655 84.855 21.975 85.405 ;
		RECT	0.32 85.955 21.655 86.735 ;
		RECT	0 85.955 0.32 86.735 ;
		RECT	21.655 85.955 21.975 86.735 ;
		RECT	0.32 87.735 21.655 88.285 ;
		RECT	0 87.735 0.32 88.285 ;
		RECT	21.655 87.735 21.975 88.285 ;
		RECT	0.32 88.835 21.655 89.615 ;
		RECT	0 88.835 0.32 89.615 ;
		RECT	21.655 88.835 21.975 89.615 ;
		RECT	0.32 90.615 21.655 91.165 ;
		RECT	0 90.615 0.32 91.165 ;
		RECT	21.655 90.615 21.975 91.165 ;
		RECT	0.32 91.715 21.655 92.495 ;
		RECT	0 91.715 0.32 92.495 ;
		RECT	21.655 91.715 21.975 92.495 ;
		RECT	0.32 93.495 21.655 94.045 ;
		RECT	0 93.495 0.32 94.045 ;
		RECT	21.655 93.495 21.975 94.045 ;
		RECT	0.32 94.595 21.655 95.375 ;
		RECT	0 94.595 0.32 95.375 ;
		RECT	21.655 94.595 21.975 95.375 ;
		RECT	0.32 96.375 21.655 96.925 ;
		RECT	0 96.375 0.32 96.925 ;
		RECT	21.655 96.375 21.975 96.925 ;
		RECT	0.32 97.475 21.655 98.255 ;
		RECT	0 97.475 0.32 98.255 ;
		RECT	21.655 97.475 21.975 98.255 ;
		RECT	0.32 99.255 21.655 99.805 ;
		RECT	0 99.255 0.32 99.805 ;
		RECT	21.655 99.255 21.975 99.805 ;
		RECT	0.32 100.355 21.655 101.135 ;
		RECT	0 100.355 0.32 101.135 ;
		RECT	21.655 100.355 21.975 101.135 ;
		RECT	0.32 102.135 21.655 102.685 ;
		RECT	0 102.135 0.32 102.685 ;
		RECT	21.655 102.135 21.975 102.685 ;
		RECT	0.32 103.235 21.655 104.015 ;
		RECT	0 103.235 0.32 104.015 ;
		RECT	21.655 103.235 21.975 104.015 ;
		RECT	0.32 105.015 21.655 105.565 ;
		RECT	0 105.015 0.32 105.565 ;
		RECT	21.655 105.015 21.975 105.565 ;
		RECT	0.32 106.115 21.655 106.895 ;
		RECT	0 106.115 0.32 106.895 ;
		RECT	21.655 106.115 21.975 106.895 ;
		RECT	0.32 107.895 21.655 108.445 ;
		RECT	0 107.895 0.32 108.445 ;
		RECT	21.655 107.895 21.975 108.445 ;
		RECT	0.32 108.995 21.655 109.775 ;
		RECT	0 108.995 0.32 109.775 ;
		RECT	21.655 108.995 21.975 109.775 ;
		RECT	0.32 110.775 21.655 111.325 ;
		RECT	0 110.775 0.32 111.325 ;
		RECT	21.655 110.775 21.975 111.325 ;
		RECT	0.32 111.875 21.655 112.655 ;
		RECT	0 111.875 0.32 112.655 ;
		RECT	21.655 111.875 21.975 112.655 ;
		RECT	0.32 113.655 21.655 114.205 ;
		RECT	0 113.655 0.32 114.205 ;
		RECT	21.655 113.655 21.975 114.205 ;
		RECT	0.32 114.755 21.655 115.535 ;
		RECT	0 114.755 0.32 115.535 ;
		RECT	21.655 114.755 21.975 115.535 ;
		RECT	0.32 116.535 21.655 117.085 ;
		RECT	0 116.535 0.32 117.085 ;
		RECT	21.655 116.535 21.975 117.085 ;
		RECT	0.32 117.635 21.655 118.415 ;
		RECT	0 117.635 0.32 118.415 ;
		RECT	21.655 117.635 21.975 118.415 ;
		RECT	0.32 119.415 21.655 119.965 ;
		RECT	0 119.415 0.32 119.965 ;
		RECT	21.655 119.415 21.975 119.965 ;
		RECT	0.32 120.515 21.655 121.295 ;
		RECT	0 120.515 0.32 121.295 ;
		RECT	21.655 120.515 21.975 121.295 ;
		RECT	0.32 122.295 21.655 122.845 ;
		RECT	0 122.295 0.32 122.845 ;
		RECT	21.655 122.295 21.975 122.845 ;
		RECT	0.32 123.395 21.655 124.175 ;
		RECT	0 123.395 0.32 124.175 ;
		RECT	21.655 123.395 21.975 124.175 ;
		RECT	0.32 125.175 21.655 125.725 ;
		RECT	0 125.175 0.32 125.725 ;
		RECT	21.655 125.175 21.975 125.725 ;
		RECT	0.32 126.275 21.655 127.055 ;
		RECT	0 126.275 0.32 127.055 ;
		RECT	21.655 126.275 21.975 127.055 ;
		RECT	0.32 128.055 21.655 128.605 ;
		RECT	0 128.055 0.32 128.605 ;
		RECT	21.655 128.055 21.975 128.605 ;
		RECT	0.32 129.155 21.655 129.935 ;
		RECT	0 129.155 0.32 129.935 ;
		RECT	21.655 129.155 21.975 129.935 ;
		RECT	0.32 130.935 21.655 131.485 ;
		RECT	0 130.935 0.32 131.485 ;
		RECT	21.655 130.935 21.975 131.485 ;
		RECT	0.32 132.035 21.655 132.815 ;
		RECT	0 132.035 0.32 132.815 ;
		RECT	21.655 132.035 21.975 132.815 ;
		RECT	0.32 133.815 21.655 134.365 ;
		RECT	0 133.815 0.32 134.365 ;
		RECT	21.655 133.815 21.975 134.365 ;
		RECT	0.32 134.915 21.655 135.695 ;
		RECT	0 134.915 0.32 135.695 ;
		RECT	21.655 134.915 21.975 135.695 ;
		RECT	0.32 136.695 21.655 137.245 ;
		RECT	0 136.695 0.32 137.245 ;
		RECT	21.655 136.695 21.975 137.245 ;
		RECT	0.32 137.795 21.655 138.575 ;
		RECT	0 137.795 0.32 138.575 ;
		RECT	21.655 137.795 21.975 138.575 ;
		RECT	0.32 139.575 21.655 140.125 ;
		RECT	0 139.575 0.32 140.125 ;
		RECT	21.655 139.575 21.975 140.125 ;
		RECT	0.32 140.675 21.655 141.455 ;
		RECT	0 140.675 0.32 141.455 ;
		RECT	21.655 140.675 21.975 141.455 ;
		RECT	0.32 142.455 21.655 143.005 ;
		RECT	0 142.455 0.32 143.005 ;
		RECT	21.655 142.455 21.975 143.005 ;
		RECT	0.32 143.555 21.655 144.335 ;
		RECT	0 143.555 0.32 144.335 ;
		RECT	21.655 143.555 21.975 144.335 ;
		RECT	0.32 145.335 21.655 145.885 ;
		RECT	0 145.335 0.32 145.885 ;
		RECT	21.655 145.335 21.975 145.885 ;
		RECT	0.32 146.435 21.655 147.215 ;
		RECT	0 146.435 0.32 147.215 ;
		RECT	21.655 146.435 21.975 147.215 ;
		RECT	0.32 148.215 21.655 148.765 ;
		RECT	0 148.215 0.32 148.765 ;
		RECT	21.655 148.215 21.975 148.765 ;
		RECT	0.32 149.315 21.655 150.095 ;
		RECT	0 149.315 0.32 150.095 ;
		RECT	21.655 149.315 21.975 150.095 ;
		RECT	0.32 151.095 21.655 151.645 ;
		RECT	0 151.095 0.32 151.645 ;
		RECT	21.655 151.095 21.975 151.645 ;
		RECT	0.32 152.195 21.655 152.975 ;
		RECT	0 152.195 0.32 152.975 ;
		RECT	21.655 152.195 21.975 152.975 ;
		RECT	0.32 153.975 21.655 154.525 ;
		RECT	0 153.975 0.32 154.525 ;
		RECT	21.655 153.975 21.975 154.525 ;
		RECT	0.32 155.075 21.655 155.855 ;
		RECT	0 155.075 0.32 155.855 ;
		RECT	21.655 155.075 21.975 155.855 ;
		RECT	0.32 156.855 21.655 157.405 ;
		RECT	0 156.855 0.32 157.405 ;
		RECT	21.655 156.855 21.975 157.405 ;
		RECT	0.32 157.955 21.655 158.735 ;
		RECT	0 157.955 0.32 158.735 ;
		RECT	21.655 157.955 21.975 158.735 ;
		RECT	0.32 159.735 21.655 160.285 ;
		RECT	0 159.735 0.32 160.285 ;
		RECT	21.655 159.735 21.975 160.285 ;
		RECT	0.32 160.835 21.655 161.615 ;
		RECT	0 160.835 0.32 161.615 ;
		RECT	21.655 160.835 21.975 161.615 ;
		RECT	0.32 162.615 21.655 163.165 ;
		RECT	0 162.615 0.32 163.165 ;
		RECT	21.655 162.615 21.975 163.165 ;
		RECT	0.32 163.715 21.655 164.495 ;
		RECT	0 163.715 0.32 164.495 ;
		RECT	21.655 163.715 21.975 164.495 ;
		RECT	0.32 165.495 21.655 166.045 ;
		RECT	0 165.495 0.32 166.045 ;
		RECT	21.655 165.495 21.975 166.045 ;
		RECT	0.32 166.595 21.655 167.375 ;
		RECT	0 166.595 0.32 167.375 ;
		RECT	21.655 166.595 21.975 167.375 ;
		RECT	0.32 168.375 21.655 168.925 ;
		RECT	0 168.375 0.32 168.925 ;
		RECT	21.655 168.375 21.975 168.925 ;
		RECT	0.32 169.475 21.655 170.255 ;
		RECT	0 169.475 0.32 170.255 ;
		RECT	21.655 169.475 21.975 170.255 ;
		RECT	0.32 171.255 21.655 171.805 ;
		RECT	0 171.255 0.32 171.805 ;
		RECT	21.655 171.255 21.975 171.805 ;
		RECT	0.32 172.355 21.655 173.135 ;
		RECT	0 172.355 0.32 173.135 ;
		RECT	21.655 172.355 21.975 173.135 ;
		RECT	0.32 174.135 21.655 174.685 ;
		RECT	0 174.135 0.32 174.685 ;
		RECT	21.655 174.135 21.975 174.685 ;
		RECT	0.32 175.235 21.655 176.015 ;
		RECT	0 175.235 0.32 176.015 ;
		RECT	21.655 175.235 21.975 176.015 ;
		RECT	0.32 177.015 21.655 177.565 ;
		RECT	0 177.015 0.32 177.565 ;
		RECT	21.655 177.015 21.975 177.565 ;
		RECT	0.32 178.115 21.655 178.895 ;
		RECT	0 178.115 0.32 178.895 ;
		RECT	21.655 178.115 21.975 178.895 ;
		RECT	0.32 179.895 21.655 180.445 ;
		RECT	0 179.895 0.32 180.445 ;
		RECT	21.655 179.895 21.975 180.445 ;
		RECT	0.32 180.995 21.655 181.775 ;
		RECT	0 180.995 0.32 181.775 ;
		RECT	21.655 180.995 21.975 181.775 ;
		RECT	0.32 182.775 21.655 183.325 ;
		RECT	0 182.775 0.32 183.325 ;
		RECT	21.655 182.775 21.975 183.325 ;
		RECT	0.32 183.875 21.655 184.655 ;
		RECT	0 183.875 0.32 184.655 ;
		RECT	21.655 183.875 21.975 184.655 ;
		RECT	0.32 185.195 21.655 186.555 ;
		RECT	0 185.195 0.32 186.555 ;
		RECT	21.655 185.195 21.975 186.555 ;
		RECT	0.32 187.325 21.655 187.835 ;
		RECT	0 187.325 0.32 187.835 ;
		RECT	21.655 187.325 21.975 187.835 ;
		RECT	0.32 188.225 21.655 188.325 ;
		RECT	0 188.225 0.32 188.325 ;
		RECT	21.655 188.225 21.975 188.325 ;
		RECT	0.32 188.715 21.655 188.815 ;
		RECT	0 188.715 0.32 188.815 ;
		RECT	21.655 188.715 21.975 188.815 ;
		RECT	0.32 189.205 21.655 190.33 ;
		RECT	0 189.205 0.32 190.33 ;
		RECT	21.655 189.205 21.975 190.33 ;
		RECT	0.32 190.72 21.655 190.785 ;
		RECT	0 190.72 0.32 190.785 ;
		RECT	21.655 190.72 21.975 190.785 ;
		RECT	0.32 191.175 21.655 191.28 ;
		RECT	0 191.175 0.32 191.28 ;
		RECT	21.655 191.175 21.975 191.28 ;
		RECT	0.32 191.67 21.655 191.77 ;
		RECT	0 191.67 0.32 191.77 ;
		RECT	21.655 191.67 21.975 191.77 ;
		RECT	0.32 192.16 21.655 192.26 ;
		RECT	0 192.16 0.32 192.26 ;
		RECT	21.655 192.16 21.975 192.26 ;
		RECT	0.32 192.65 21.655 193.245 ;
		RECT	0 192.65 0.32 193.245 ;
		RECT	21.655 192.65 21.975 193.245 ;
		RECT	0.32 193.635 21.655 194.23 ;
		RECT	0 193.635 0.32 194.23 ;
		RECT	21.655 193.635 21.975 194.23 ;
		RECT	0.32 194.62 21.655 194.725 ;
		RECT	0 194.62 0.32 194.725 ;
		RECT	21.655 194.62 21.975 194.725 ;
		RECT	0.32 195.115 21.655 195.215 ;
		RECT	0 195.115 0.32 195.215 ;
		RECT	21.655 195.115 21.975 195.215 ;
		RECT	0.32 195.605 21.655 195.705 ;
		RECT	0 195.605 0.32 195.705 ;
		RECT	21.655 195.605 21.975 195.705 ;
		RECT	0.32 196.095 21.655 196.2 ;
		RECT	0 196.095 0.32 196.2 ;
		RECT	21.655 196.095 21.975 196.2 ;
		RECT	0.32 196.59 21.655 196.69 ;
		RECT	0 196.59 0.32 196.69 ;
		RECT	21.655 196.59 21.975 196.69 ;
		RECT	0.32 197.08 21.655 197.18 ;
		RECT	0 197.08 0.32 197.18 ;
		RECT	21.655 197.08 21.975 197.18 ;
		RECT	0.32 197.57 21.655 198.165 ;
		RECT	0 197.57 0.32 198.165 ;
		RECT	21.655 197.57 21.975 198.165 ;
		RECT	0.32 198.555 21.655 198.66 ;
		RECT	0 198.555 0.32 198.66 ;
		RECT	21.655 198.555 21.975 198.66 ;
		RECT	0.32 199.05 21.655 199.15 ;
		RECT	0 199.05 0.32 199.15 ;
		RECT	21.655 199.05 21.975 199.15 ;
		RECT	0.32 199.54 21.655 199.63 ;
		RECT	0 199.54 0.32 199.63 ;
		RECT	21.655 199.54 21.975 199.63 ;
		RECT	0.32 200.04 21.655 200.135 ;
		RECT	0 200.04 0.32 200.135 ;
		RECT	21.655 200.04 21.975 200.135 ;
		RECT	0.32 200.525 21.655 200.625 ;
		RECT	0 200.525 0.32 200.625 ;
		RECT	21.655 200.525 21.975 200.625 ;
		RECT	0.32 201.015 21.655 201.12 ;
		RECT	0 201.015 0.32 201.12 ;
		RECT	21.655 201.015 21.975 201.12 ;
		RECT	0.32 201.51 21.655 202.6 ;
		RECT	0 201.51 0.32 202.6 ;
		RECT	21.655 201.51 21.975 202.6 ;
		RECT	0.32 202.99 21.655 203.085 ;
		RECT	0 202.99 0.32 203.085 ;
		RECT	21.655 202.99 21.975 203.085 ;
		RECT	0.32 203.475 21.655 203.58 ;
		RECT	0 203.475 0.32 203.58 ;
		RECT	21.655 203.475 21.975 203.58 ;
		RECT	0.32 203.97 21.655 205.055 ;
		RECT	0 203.97 0.32 205.055 ;
		RECT	21.655 203.97 21.975 205.055 ;
		RECT	0.32 205.445 21.655 206.04 ;
		RECT	0 205.445 0.32 206.04 ;
		RECT	21.655 205.445 21.975 206.04 ;
		RECT	0.32 206.43 21.655 206.53 ;
		RECT	0 206.43 0.32 206.53 ;
		RECT	21.655 206.43 21.975 206.53 ;
		RECT	0.32 206.92 21.655 207.02 ;
		RECT	0 206.92 0.32 207.02 ;
		RECT	21.655 206.92 21.975 207.02 ;
		RECT	0.32 207.41 21.655 207.515 ;
		RECT	0 207.41 0.32 207.515 ;
		RECT	21.655 207.41 21.975 207.515 ;
		RECT	0.32 207.905 21.655 208.005 ;
		RECT	0 207.905 0.32 208.005 ;
		RECT	21.655 207.905 21.975 208.005 ;
		RECT	0.32 208.395 21.655 208.5 ;
		RECT	0 208.395 0.32 208.5 ;
		RECT	21.655 208.395 21.975 208.5 ;
		RECT	0.32 208.89 21.655 209.48 ;
		RECT	0 208.89 0.32 209.48 ;
		RECT	21.655 208.89 21.975 209.48 ;
		RECT	0.32 209.87 21.655 210.955 ;
		RECT	0 209.87 0.32 210.955 ;
		RECT	21.655 209.87 21.975 210.955 ;
		RECT	0.32 211.345 21.655 211.45 ;
		RECT	0 211.345 0.32 211.45 ;
		RECT	21.655 211.345 21.975 211.45 ;
		RECT	0.32 211.84 21.655 211.945 ;
		RECT	0 211.84 0.32 211.945 ;
		RECT	21.655 211.84 21.975 211.945 ;
		RECT	0.32 212.335 21.655 213.42 ;
		RECT	0 212.335 0.32 213.42 ;
		RECT	21.655 212.335 21.975 213.42 ;
		RECT	0.32 213.81 21.655 213.91 ;
		RECT	0 213.81 0.32 213.91 ;
		RECT	21.655 213.81 21.975 213.91 ;
		RECT	0.32 214.3 21.655 214.405 ;
		RECT	0 214.3 0.32 214.405 ;
		RECT	21.655 214.3 21.975 214.405 ;
		RECT	0.32 214.795 21.655 214.885 ;
		RECT	0 214.795 0.32 214.885 ;
		RECT	21.655 214.795 21.975 214.885 ;
		RECT	0.32 215.295 21.655 215.385 ;
		RECT	0 215.295 0.32 215.385 ;
		RECT	21.655 215.295 21.975 215.385 ;
		RECT	0.32 215.775 21.655 215.88 ;
		RECT	0 215.775 0.32 215.88 ;
		RECT	21.655 215.775 21.975 215.88 ;
		RECT	0.32 216.27 21.655 216.37 ;
		RECT	0 216.27 0.32 216.37 ;
		RECT	21.655 216.27 21.975 216.37 ;
		RECT	0.32 216.76 21.655 217.355 ;
		RECT	0 216.76 0.32 217.355 ;
		RECT	21.655 216.76 21.975 217.355 ;
		RECT	0.32 217.745 21.655 217.845 ;
		RECT	0 217.745 0.32 217.845 ;
		RECT	21.655 217.745 21.975 217.845 ;
		RECT	0.32 218.235 21.655 218.34 ;
		RECT	0 218.235 0.32 218.34 ;
		RECT	21.655 218.235 21.975 218.34 ;
		RECT	0.32 218.73 21.655 218.83 ;
		RECT	0 218.73 0.32 218.83 ;
		RECT	21.655 218.73 21.975 218.83 ;
		RECT	0.32 219.22 21.655 219.325 ;
		RECT	0 219.22 0.32 219.325 ;
		RECT	21.655 219.22 21.975 219.325 ;
		RECT	0.32 219.715 21.655 219.815 ;
		RECT	0 219.715 0.32 219.815 ;
		RECT	21.655 219.715 21.975 219.815 ;
		RECT	0.32 220.205 21.655 220.305 ;
		RECT	0 220.205 0.32 220.305 ;
		RECT	21.655 220.205 21.975 220.305 ;
		RECT	0.32 220.695 21.655 221.29 ;
		RECT	0 220.695 0.32 221.29 ;
		RECT	21.655 220.695 21.975 221.29 ;
		RECT	0.32 221.68 21.655 222.275 ;
		RECT	0 221.68 0.32 222.275 ;
		RECT	21.655 221.68 21.975 222.275 ;
		RECT	0.32 222.665 21.655 222.755 ;
		RECT	0 222.665 0.32 222.755 ;
		RECT	21.655 222.665 21.975 222.755 ;
		RECT	0.32 223.165 21.655 223.225 ;
		RECT	0 223.165 0.32 223.225 ;
		RECT	21.655 223.165 21.975 223.225 ;
		RECT	0.32 223.615 21.655 223.75 ;
		RECT	0 223.615 0.32 223.75 ;
		RECT	21.655 223.615 21.975 223.75 ;
		RECT	0.32 224.14 21.655 224.21 ;
		RECT	0 224.14 0.32 224.21 ;
		RECT	21.655 224.14 21.975 224.21 ;
		RECT	0.32 224.6 21.655 225.72 ;
		RECT	0 224.6 0.32 225.72 ;
		RECT	21.655 224.6 21.975 225.72 ;
		RECT	0.32 226.11 21.655 226.21 ;
		RECT	0 226.11 0.32 226.21 ;
		RECT	21.655 226.11 21.975 226.21 ;
		RECT	0.32 226.6 21.655 226.705 ;
		RECT	0 226.6 0.32 226.705 ;
		RECT	21.655 226.6 21.975 226.705 ;
		RECT	0.32 227.095 21.655 227.535 ;
		RECT	0 227.095 0.32 227.535 ;
		RECT	21.655 227.095 21.975 227.535 ;
		RECT	0.32 228.305 21.655 229.665 ;
		RECT	0 228.305 0.32 229.665 ;
		RECT	21.655 228.305 21.975 229.665 ;
		RECT	0.32 230.205 21.655 230.985 ;
		RECT	0 230.205 0.32 230.985 ;
		RECT	21.655 230.205 21.975 230.985 ;
		RECT	0.32 231.535 21.655 232.085 ;
		RECT	0 231.535 0.32 232.085 ;
		RECT	21.655 231.535 21.975 232.085 ;
		RECT	0.32 233.085 21.655 233.865 ;
		RECT	0 233.085 0.32 233.865 ;
		RECT	21.655 233.085 21.975 233.865 ;
		RECT	0.32 234.415 21.655 234.965 ;
		RECT	0 234.415 0.32 234.965 ;
		RECT	21.655 234.415 21.975 234.965 ;
		RECT	0.32 235.965 21.655 236.745 ;
		RECT	0 235.965 0.32 236.745 ;
		RECT	21.655 235.965 21.975 236.745 ;
		RECT	0.32 237.295 21.655 237.845 ;
		RECT	0 237.295 0.32 237.845 ;
		RECT	21.655 237.295 21.975 237.845 ;
		RECT	0.32 238.845 21.655 239.625 ;
		RECT	0 238.845 0.32 239.625 ;
		RECT	21.655 238.845 21.975 239.625 ;
		RECT	0.32 240.175 21.655 240.725 ;
		RECT	0 240.175 0.32 240.725 ;
		RECT	21.655 240.175 21.975 240.725 ;
		RECT	0.32 241.725 21.655 242.505 ;
		RECT	0 241.725 0.32 242.505 ;
		RECT	21.655 241.725 21.975 242.505 ;
		RECT	0.32 243.055 21.655 243.605 ;
		RECT	0 243.055 0.32 243.605 ;
		RECT	21.655 243.055 21.975 243.605 ;
		RECT	0.32 244.605 21.655 245.385 ;
		RECT	0 244.605 0.32 245.385 ;
		RECT	21.655 244.605 21.975 245.385 ;
		RECT	0.32 245.935 21.655 246.485 ;
		RECT	0 245.935 0.32 246.485 ;
		RECT	21.655 245.935 21.975 246.485 ;
		RECT	0.32 247.485 21.655 248.265 ;
		RECT	0 247.485 0.32 248.265 ;
		RECT	21.655 247.485 21.975 248.265 ;
		RECT	0.32 248.815 21.655 249.365 ;
		RECT	0 248.815 0.32 249.365 ;
		RECT	21.655 248.815 21.975 249.365 ;
		RECT	0.32 250.365 21.655 251.145 ;
		RECT	0 250.365 0.32 251.145 ;
		RECT	21.655 250.365 21.975 251.145 ;
		RECT	0.32 251.695 21.655 252.245 ;
		RECT	0 251.695 0.32 252.245 ;
		RECT	21.655 251.695 21.975 252.245 ;
		RECT	0.32 253.245 21.655 254.025 ;
		RECT	0 253.245 0.32 254.025 ;
		RECT	21.655 253.245 21.975 254.025 ;
		RECT	0.32 254.575 21.655 255.125 ;
		RECT	0 254.575 0.32 255.125 ;
		RECT	21.655 254.575 21.975 255.125 ;
		RECT	0.32 256.125 21.655 256.905 ;
		RECT	0 256.125 0.32 256.905 ;
		RECT	21.655 256.125 21.975 256.905 ;
		RECT	0.32 257.455 21.655 258.005 ;
		RECT	0 257.455 0.32 258.005 ;
		RECT	21.655 257.455 21.975 258.005 ;
		RECT	0.32 259.005 21.655 259.785 ;
		RECT	0 259.005 0.32 259.785 ;
		RECT	21.655 259.005 21.975 259.785 ;
		RECT	0.32 260.335 21.655 260.885 ;
		RECT	0 260.335 0.32 260.885 ;
		RECT	21.655 260.335 21.975 260.885 ;
		RECT	0.32 261.885 21.655 262.665 ;
		RECT	0 261.885 0.32 262.665 ;
		RECT	21.655 261.885 21.975 262.665 ;
		RECT	0.32 263.215 21.655 263.765 ;
		RECT	0 263.215 0.32 263.765 ;
		RECT	21.655 263.215 21.975 263.765 ;
		RECT	0.32 264.765 21.655 265.545 ;
		RECT	0 264.765 0.32 265.545 ;
		RECT	21.655 264.765 21.975 265.545 ;
		RECT	0.32 266.095 21.655 266.645 ;
		RECT	0 266.095 0.32 266.645 ;
		RECT	21.655 266.095 21.975 266.645 ;
		RECT	0.32 267.645 21.655 268.425 ;
		RECT	0 267.645 0.32 268.425 ;
		RECT	21.655 267.645 21.975 268.425 ;
		RECT	0.32 268.975 21.655 269.525 ;
		RECT	0 268.975 0.32 269.525 ;
		RECT	21.655 268.975 21.975 269.525 ;
		RECT	0.32 270.525 21.655 271.305 ;
		RECT	0 270.525 0.32 271.305 ;
		RECT	21.655 270.525 21.975 271.305 ;
		RECT	0.32 271.855 21.655 272.405 ;
		RECT	0 271.855 0.32 272.405 ;
		RECT	21.655 271.855 21.975 272.405 ;
		RECT	0.32 273.405 21.655 274.185 ;
		RECT	0 273.405 0.32 274.185 ;
		RECT	21.655 273.405 21.975 274.185 ;
		RECT	0.32 274.735 21.655 275.285 ;
		RECT	0 274.735 0.32 275.285 ;
		RECT	21.655 274.735 21.975 275.285 ;
		RECT	0.32 276.285 21.655 277.065 ;
		RECT	0 276.285 0.32 277.065 ;
		RECT	21.655 276.285 21.975 277.065 ;
		RECT	0.32 277.615 21.655 278.165 ;
		RECT	0 277.615 0.32 278.165 ;
		RECT	21.655 277.615 21.975 278.165 ;
		RECT	0.32 279.165 21.655 279.945 ;
		RECT	0 279.165 0.32 279.945 ;
		RECT	21.655 279.165 21.975 279.945 ;
		RECT	0.32 280.495 21.655 281.045 ;
		RECT	0 280.495 0.32 281.045 ;
		RECT	21.655 280.495 21.975 281.045 ;
		RECT	0.32 282.045 21.655 282.825 ;
		RECT	0 282.045 0.32 282.825 ;
		RECT	21.655 282.045 21.975 282.825 ;
		RECT	0.32 283.375 21.655 283.925 ;
		RECT	0 283.375 0.32 283.925 ;
		RECT	21.655 283.375 21.975 283.925 ;
		RECT	0.32 284.925 21.655 285.705 ;
		RECT	0 284.925 0.32 285.705 ;
		RECT	21.655 284.925 21.975 285.705 ;
		RECT	0.32 286.255 21.655 286.805 ;
		RECT	0 286.255 0.32 286.805 ;
		RECT	21.655 286.255 21.975 286.805 ;
		RECT	0.32 287.805 21.655 288.585 ;
		RECT	0 287.805 0.32 288.585 ;
		RECT	21.655 287.805 21.975 288.585 ;
		RECT	0.32 289.135 21.655 289.685 ;
		RECT	0 289.135 0.32 289.685 ;
		RECT	21.655 289.135 21.975 289.685 ;
		RECT	0.32 290.685 21.655 291.465 ;
		RECT	0 290.685 0.32 291.465 ;
		RECT	21.655 290.685 21.975 291.465 ;
		RECT	0.32 292.015 21.655 292.565 ;
		RECT	0 292.015 0.32 292.565 ;
		RECT	21.655 292.015 21.975 292.565 ;
		RECT	0.32 293.565 21.655 294.345 ;
		RECT	0 293.565 0.32 294.345 ;
		RECT	21.655 293.565 21.975 294.345 ;
		RECT	0.32 294.895 21.655 295.445 ;
		RECT	0 294.895 0.32 295.445 ;
		RECT	21.655 294.895 21.975 295.445 ;
		RECT	0.32 296.445 21.655 297.225 ;
		RECT	0 296.445 0.32 297.225 ;
		RECT	21.655 296.445 21.975 297.225 ;
		RECT	0.32 297.775 21.655 298.325 ;
		RECT	0 297.775 0.32 298.325 ;
		RECT	21.655 297.775 21.975 298.325 ;
		RECT	0.32 299.325 21.655 300.105 ;
		RECT	0 299.325 0.32 300.105 ;
		RECT	21.655 299.325 21.975 300.105 ;
		RECT	0.32 300.655 21.655 301.205 ;
		RECT	0 300.655 0.32 301.205 ;
		RECT	21.655 300.655 21.975 301.205 ;
		RECT	0.32 302.205 21.655 302.985 ;
		RECT	0 302.205 0.32 302.985 ;
		RECT	21.655 302.205 21.975 302.985 ;
		RECT	0.32 303.535 21.655 304.085 ;
		RECT	0 303.535 0.32 304.085 ;
		RECT	21.655 303.535 21.975 304.085 ;
		RECT	0.32 305.085 21.655 305.865 ;
		RECT	0 305.085 0.32 305.865 ;
		RECT	21.655 305.085 21.975 305.865 ;
		RECT	0.32 306.415 21.655 306.965 ;
		RECT	0 306.415 0.32 306.965 ;
		RECT	21.655 306.415 21.975 306.965 ;
		RECT	0.32 307.965 21.655 308.745 ;
		RECT	0 307.965 0.32 308.745 ;
		RECT	21.655 307.965 21.975 308.745 ;
		RECT	0.32 309.295 21.655 309.845 ;
		RECT	0 309.295 0.32 309.845 ;
		RECT	21.655 309.295 21.975 309.845 ;
		RECT	0.32 310.845 21.655 311.625 ;
		RECT	0 310.845 0.32 311.625 ;
		RECT	21.655 310.845 21.975 311.625 ;
		RECT	0.32 312.175 21.655 312.725 ;
		RECT	0 312.175 0.32 312.725 ;
		RECT	21.655 312.175 21.975 312.725 ;
		RECT	0.32 313.725 21.655 314.505 ;
		RECT	0 313.725 0.32 314.505 ;
		RECT	21.655 313.725 21.975 314.505 ;
		RECT	0.32 315.055 21.655 315.605 ;
		RECT	0 315.055 0.32 315.605 ;
		RECT	21.655 315.055 21.975 315.605 ;
		RECT	0.32 316.605 21.655 317.385 ;
		RECT	0 316.605 0.32 317.385 ;
		RECT	21.655 316.605 21.975 317.385 ;
		RECT	0.32 317.935 21.655 318.485 ;
		RECT	0 317.935 0.32 318.485 ;
		RECT	21.655 317.935 21.975 318.485 ;
		RECT	0.32 319.485 21.655 320.265 ;
		RECT	0 319.485 0.32 320.265 ;
		RECT	21.655 319.485 21.975 320.265 ;
		RECT	0.32 320.815 21.655 321.365 ;
		RECT	0 320.815 0.32 321.365 ;
		RECT	21.655 320.815 21.975 321.365 ;
		RECT	0.32 322.365 21.655 323.145 ;
		RECT	0 322.365 0.32 323.145 ;
		RECT	21.655 322.365 21.975 323.145 ;
		RECT	0.32 323.695 21.655 324.245 ;
		RECT	0 323.695 0.32 324.245 ;
		RECT	21.655 323.695 21.975 324.245 ;
		RECT	0.32 325.245 21.655 326.025 ;
		RECT	0 325.245 0.32 326.025 ;
		RECT	21.655 325.245 21.975 326.025 ;
		RECT	0.32 326.575 21.655 327.125 ;
		RECT	0 326.575 0.32 327.125 ;
		RECT	21.655 326.575 21.975 327.125 ;
		RECT	0.32 328.125 21.655 328.905 ;
		RECT	0 328.125 0.32 328.905 ;
		RECT	21.655 328.125 21.975 328.905 ;
		RECT	0.32 329.455 21.655 330.005 ;
		RECT	0 329.455 0.32 330.005 ;
		RECT	21.655 329.455 21.975 330.005 ;
		RECT	0.32 331.005 21.655 331.785 ;
		RECT	0 331.005 0.32 331.785 ;
		RECT	21.655 331.005 21.975 331.785 ;
		RECT	0.32 332.335 21.655 332.885 ;
		RECT	0 332.335 0.32 332.885 ;
		RECT	21.655 332.335 21.975 332.885 ;
		RECT	0.32 333.885 21.655 334.665 ;
		RECT	0 333.885 0.32 334.665 ;
		RECT	21.655 333.885 21.975 334.665 ;
		RECT	0.32 335.215 21.655 335.765 ;
		RECT	0 335.215 0.32 335.765 ;
		RECT	21.655 335.215 21.975 335.765 ;
		RECT	0.32 336.765 21.655 337.545 ;
		RECT	0 336.765 0.32 337.545 ;
		RECT	21.655 336.765 21.975 337.545 ;
		RECT	0.32 338.095 21.655 338.645 ;
		RECT	0 338.095 0.32 338.645 ;
		RECT	21.655 338.095 21.975 338.645 ;
		RECT	0.32 339.645 21.655 340.425 ;
		RECT	0 339.645 0.32 340.425 ;
		RECT	21.655 339.645 21.975 340.425 ;
		RECT	0.32 340.975 21.655 341.525 ;
		RECT	0 340.975 0.32 341.525 ;
		RECT	21.655 340.975 21.975 341.525 ;
		RECT	0.32 342.525 21.655 343.305 ;
		RECT	0 342.525 0.32 343.305 ;
		RECT	21.655 342.525 21.975 343.305 ;
		RECT	0.32 343.855 21.655 344.405 ;
		RECT	0 343.855 0.32 344.405 ;
		RECT	21.655 343.855 21.975 344.405 ;
		RECT	0.32 345.405 21.655 346.185 ;
		RECT	0 345.405 0.32 346.185 ;
		RECT	21.655 345.405 21.975 346.185 ;
		RECT	0.32 346.735 21.655 347.285 ;
		RECT	0 346.735 0.32 347.285 ;
		RECT	21.655 346.735 21.975 347.285 ;
		RECT	0.32 348.285 21.655 349.065 ;
		RECT	0 348.285 0.32 349.065 ;
		RECT	21.655 348.285 21.975 349.065 ;
		RECT	0.32 349.615 21.655 350.165 ;
		RECT	0 349.615 0.32 350.165 ;
		RECT	21.655 349.615 21.975 350.165 ;
		RECT	0.32 351.165 21.655 351.945 ;
		RECT	0 351.165 0.32 351.945 ;
		RECT	21.655 351.165 21.975 351.945 ;
		RECT	0.32 352.495 21.655 353.045 ;
		RECT	0 352.495 0.32 353.045 ;
		RECT	21.655 352.495 21.975 353.045 ;
		RECT	0.32 354.045 21.655 354.825 ;
		RECT	0 354.045 0.32 354.825 ;
		RECT	21.655 354.045 21.975 354.825 ;
		RECT	0.32 355.375 21.655 355.925 ;
		RECT	0 355.375 0.32 355.925 ;
		RECT	21.655 355.375 21.975 355.925 ;
		RECT	0.32 356.925 21.655 357.705 ;
		RECT	0 356.925 0.32 357.705 ;
		RECT	21.655 356.925 21.975 357.705 ;
		RECT	0.32 358.255 21.655 358.805 ;
		RECT	0 358.255 0.32 358.805 ;
		RECT	21.655 358.255 21.975 358.805 ;
		RECT	0.32 359.805 21.655 360.585 ;
		RECT	0 359.805 0.32 360.585 ;
		RECT	21.655 359.805 21.975 360.585 ;
		RECT	0.32 361.135 21.655 361.685 ;
		RECT	0 361.135 0.32 361.685 ;
		RECT	21.655 361.135 21.975 361.685 ;
		RECT	0.32 362.685 21.655 363.465 ;
		RECT	0 362.685 0.32 363.465 ;
		RECT	21.655 362.685 21.975 363.465 ;
		RECT	0.32 364.015 21.655 364.565 ;
		RECT	0 364.015 0.32 364.565 ;
		RECT	21.655 364.015 21.975 364.565 ;
		RECT	0.32 365.565 21.655 366.345 ;
		RECT	0 365.565 0.32 366.345 ;
		RECT	21.655 365.565 21.975 366.345 ;
		RECT	0.32 366.895 21.655 367.445 ;
		RECT	0 366.895 0.32 367.445 ;
		RECT	21.655 366.895 21.975 367.445 ;
		RECT	0.32 368.445 21.655 369.225 ;
		RECT	0 368.445 0.32 369.225 ;
		RECT	21.655 368.445 21.975 369.225 ;
		RECT	0.32 369.775 21.655 370.325 ;
		RECT	0 369.775 0.32 370.325 ;
		RECT	21.655 369.775 21.975 370.325 ;
		RECT	0.32 371.325 21.655 372.105 ;
		RECT	0 371.325 0.32 372.105 ;
		RECT	21.655 371.325 21.975 372.105 ;
		RECT	0.32 372.655 21.655 373.205 ;
		RECT	0 372.655 0.32 373.205 ;
		RECT	21.655 372.655 21.975 373.205 ;
		RECT	0.32 374.205 21.655 374.985 ;
		RECT	0 374.205 0.32 374.985 ;
		RECT	21.655 374.205 21.975 374.985 ;
		RECT	0.32 375.535 21.655 376.085 ;
		RECT	0 375.535 0.32 376.085 ;
		RECT	21.655 375.535 21.975 376.085 ;
		RECT	0.32 377.085 21.655 377.865 ;
		RECT	0 377.085 0.32 377.865 ;
		RECT	21.655 377.085 21.975 377.865 ;
		RECT	0.32 378.415 21.655 378.965 ;
		RECT	0 378.415 0.32 378.965 ;
		RECT	21.655 378.415 21.975 378.965 ;
		RECT	0.32 379.965 21.655 380.745 ;
		RECT	0 379.965 0.32 380.745 ;
		RECT	21.655 379.965 21.975 380.745 ;
		RECT	0.32 381.295 21.655 381.845 ;
		RECT	0 381.295 0.32 381.845 ;
		RECT	21.655 381.295 21.975 381.845 ;
		RECT	0.32 382.845 21.655 383.625 ;
		RECT	0 382.845 0.32 383.625 ;
		RECT	21.655 382.845 21.975 383.625 ;
		RECT	0.32 384.175 21.655 384.725 ;
		RECT	0 384.175 0.32 384.725 ;
		RECT	21.655 384.175 21.975 384.725 ;
		RECT	0.32 385.725 21.655 386.505 ;
		RECT	0 385.725 0.32 386.505 ;
		RECT	21.655 385.725 21.975 386.505 ;
		RECT	0.32 387.055 21.655 387.605 ;
		RECT	0 387.055 0.32 387.605 ;
		RECT	21.655 387.055 21.975 387.605 ;
		RECT	0.32 388.605 21.655 389.385 ;
		RECT	0 388.605 0.32 389.385 ;
		RECT	21.655 388.605 21.975 389.385 ;
		RECT	0.32 389.935 21.655 390.485 ;
		RECT	0 389.935 0.32 390.485 ;
		RECT	21.655 389.935 21.975 390.485 ;
		RECT	0.32 391.485 21.655 392.265 ;
		RECT	0 391.485 0.32 392.265 ;
		RECT	21.655 391.485 21.975 392.265 ;
		RECT	0.32 392.815 21.655 393.365 ;
		RECT	0 392.815 0.32 393.365 ;
		RECT	21.655 392.815 21.975 393.365 ;
		RECT	0.32 394.365 21.655 395.145 ;
		RECT	0 394.365 0.32 395.145 ;
		RECT	21.655 394.365 21.975 395.145 ;
		RECT	0.32 395.695 21.655 396.245 ;
		RECT	0 395.695 0.32 396.245 ;
		RECT	21.655 395.695 21.975 396.245 ;
		RECT	0.32 397.245 21.655 398.025 ;
		RECT	0 397.245 0.32 398.025 ;
		RECT	21.655 397.245 21.975 398.025 ;
		RECT	0.32 398.575 21.655 399.125 ;
		RECT	0 398.575 0.32 399.125 ;
		RECT	21.655 398.575 21.975 399.125 ;
		RECT	0.32 400.125 21.655 400.905 ;
		RECT	0 400.125 0.32 400.905 ;
		RECT	21.655 400.125 21.975 400.905 ;
		RECT	0.32 401.455 21.655 402.005 ;
		RECT	0 401.455 0.32 402.005 ;
		RECT	21.655 401.455 21.975 402.005 ;
		RECT	0.32 403.005 21.655 403.785 ;
		RECT	0 403.005 0.32 403.785 ;
		RECT	21.655 403.005 21.975 403.785 ;
		RECT	0.32 404.335 21.655 404.885 ;
		RECT	0 404.335 0.32 404.885 ;
		RECT	21.655 404.335 21.975 404.885 ;
		RECT	0.32 405.885 21.655 406.665 ;
		RECT	0 405.885 0.32 406.665 ;
		RECT	21.655 405.885 21.975 406.665 ;
		RECT	0.32 407.215 21.655 407.765 ;
		RECT	0 407.215 0.32 407.765 ;
		RECT	21.655 407.215 21.975 407.765 ;
		RECT	0.32 408.765 21.655 409.545 ;
		RECT	0 408.765 0.32 409.545 ;
		RECT	21.655 408.765 21.975 409.545 ;
		RECT	0.32 410.095 21.655 410.645 ;
		RECT	0 410.095 0.32 410.645 ;
		RECT	21.655 410.095 21.975 410.645 ;
		RECT	0.32 411.645 21.655 412.425 ;
		RECT	0 411.645 0.32 412.425 ;
		RECT	21.655 411.645 21.975 412.425 ;
		RECT	0.32 412.975 21.655 413.525 ;
		RECT	0 412.975 0.32 413.525 ;
		RECT	21.655 412.975 21.975 413.525 ;
		RECT	0.32 414.755 21.655 414.86 ;
		RECT	0 414.755 0.32 414.86 ;
		RECT	21.655 414.755 21.975 414.86 ;
		LAYER	VIA1 DESIGNRULEWIDTH 0.07 ;
		RECT	0 0 21.975 414.86 ;
		LAYER	VIA2 DESIGNRULEWIDTH 0.07 ;
		RECT	0 0 21.975 414.86 ;
		LAYER	VIA3 DESIGNRULEWIDTH 0.07 ;
		RECT	0.435 186.415 0.485 186.545 ;
		RECT	0.435 187.58 0.485 187.71 ;
		RECT	0.435 189.445 0.485 189.575 ;
		RECT	0.435 189.915 0.485 190.045 ;
		RECT	0.435 193.87 0.485 194 ;
		RECT	0.435 197.805 0.485 197.935 ;
		RECT	0.435 201.74 0.485 201.87 ;
		RECT	0.435 204.865 0.485 204.995 ;
		RECT	0.435 205.675 0.485 205.805 ;
		RECT	0.435 209.12 0.485 209.25 ;
		RECT	0.435 209.93 0.485 210.06 ;
		RECT	0.435 213.055 0.485 213.185 ;
		RECT	0.435 216.995 0.485 217.125 ;
		RECT	0.435 220.93 0.485 221.06 ;
		RECT	0.435 224.88 0.485 225.01 ;
		RECT	0.435 225.355 0.485 225.485 ;
		RECT	0.435 227.145 0.485 227.275 ;
		RECT	0.435 228.315 0.485 228.445 ;
		RECT	0.435 186.875 0.485 187.005 ;
		RECT	0.435 192.885 0.485 193.015 ;
		RECT	0.435 221.915 0.485 222.045 ;
		RECT	0.435 227.855 0.485 227.985 ;
		RECT	1.625 186.415 1.675 186.545 ;
		RECT	1.92 186.415 1.97 186.545 ;
		RECT	2.4 186.415 2.45 186.545 ;
		RECT	2.55 186.415 2.6 186.545 ;
		RECT	3.79 186.415 3.84 186.545 ;
		RECT	4.055 186.415 4.105 186.545 ;
		RECT	5.05 186.415 5.1 186.545 ;
		RECT	5.575 186.415 5.625 186.545 ;
		RECT	6.76 186.415 6.81 186.545 ;
		RECT	8.04 186.415 8.09 186.545 ;
		RECT	9.855 186.415 9.905 186.545 ;
		RECT	10.26 186.415 10.31 186.545 ;
		RECT	11.565 186.415 11.615 186.545 ;
		RECT	0.62 186.645 0.67 186.775 ;
		RECT	1.16 186.645 1.21 186.775 ;
		RECT	4.19 186.645 4.24 186.775 ;
		RECT	7.73 186.645 7.78 186.775 ;
		RECT	14.68 186.645 14.73 186.775 ;
		RECT	2.72 186.875 2.77 187.005 ;
		RECT	9.1 186.875 9.15 187.005 ;
		RECT	10.81 186.875 10.86 187.005 ;
		RECT	14.34 187.105 14.39 187.235 ;
		RECT	2.4 187.58 2.45 187.71 ;
		RECT	2.55 187.58 2.6 187.71 ;
		RECT	3.79 187.58 3.84 187.71 ;
		RECT	4.055 187.58 4.105 187.71 ;
		RECT	5.575 187.58 5.625 187.71 ;
		RECT	6.76 187.58 6.81 187.71 ;
		RECT	8.04 187.58 8.09 187.71 ;
		RECT	10.26 187.58 10.31 187.71 ;
		RECT	11.565 187.58 11.615 187.71 ;
		RECT	1.585 187.62 1.715 187.67 ;
		RECT	1.88 187.62 2.01 187.67 ;
		RECT	5.01 187.62 5.14 187.67 ;
		RECT	9.815 187.62 9.945 187.67 ;
		RECT	2.11 187.965 2.16 188.095 ;
		RECT	5.41 187.965 5.46 188.095 ;
		RECT	6.44 187.965 6.49 188.095 ;
		RECT	9.495 187.965 9.545 188.095 ;
		RECT	13.33 187.965 13.38 188.095 ;
		RECT	14.87 187.965 14.92 188.095 ;
		RECT	15.065 187.965 15.115 188.095 ;
		RECT	3.56 188.005 3.69 188.055 ;
		RECT	0.9 188.455 0.95 188.585 ;
		RECT	1.44 188.455 1.49 188.585 ;
		RECT	3.025 188.455 3.075 188.585 ;
		RECT	3.155 188.455 3.205 188.585 ;
		RECT	6.605 188.455 6.655 188.585 ;
		RECT	7.265 188.455 7.315 188.585 ;
		RECT	12.095 188.455 12.145 188.585 ;
		RECT	12.355 188.455 12.405 188.585 ;
		RECT	13.06 188.455 13.11 188.585 ;
		RECT	14.545 188.455 14.595 188.585 ;
		RECT	4.34 188.495 4.47 188.545 ;
		RECT	6.175 188.495 6.305 188.545 ;
		RECT	8.85 188.495 8.98 188.545 ;
		RECT	9.27 188.495 9.4 188.545 ;
		RECT	12.225 188.74 12.275 188.79 ;
		RECT	13.195 188.74 13.245 188.79 ;
		RECT	2.11 188.945 2.16 189.075 ;
		RECT	5.41 188.945 5.46 189.075 ;
		RECT	6.44 188.945 6.49 189.075 ;
		RECT	9.495 188.945 9.545 189.075 ;
		RECT	13.33 188.945 13.38 189.075 ;
		RECT	14.875 188.945 14.925 189.075 ;
		RECT	15.07 188.945 15.12 189.075 ;
		RECT	3.56 188.985 3.69 189.035 ;
		RECT	1.585 189.42 1.715 189.47 ;
		RECT	1.88 189.42 2.01 189.47 ;
		RECT	5.01 189.42 5.14 189.47 ;
		RECT	9.815 189.42 9.945 189.47 ;
		RECT	14.215 189.44 14.265 189.57 ;
		RECT	2.4 189.445 2.45 189.575 ;
		RECT	2.55 189.445 2.6 189.575 ;
		RECT	3.79 189.445 3.84 189.575 ;
		RECT	4.055 189.445 4.105 189.575 ;
		RECT	5.575 189.445 5.625 189.575 ;
		RECT	6.76 189.445 6.81 189.575 ;
		RECT	8.04 189.445 8.09 189.575 ;
		RECT	10.26 189.445 10.31 189.575 ;
		RECT	11.565 189.445 11.615 189.575 ;
		RECT	1.585 189.55 1.715 189.6 ;
		RECT	1.88 189.55 2.01 189.6 ;
		RECT	5.01 189.55 5.14 189.6 ;
		RECT	9.815 189.55 9.945 189.6 ;
		RECT	12.225 189.72 12.275 189.77 ;
		RECT	13.195 189.72 13.245 189.77 ;
		RECT	2.4 189.915 2.45 190.045 ;
		RECT	2.55 189.915 2.6 190.045 ;
		RECT	3.79 189.915 3.84 190.045 ;
		RECT	4.055 189.915 4.105 190.045 ;
		RECT	5.575 189.915 5.625 190.045 ;
		RECT	6.76 189.915 6.81 190.045 ;
		RECT	8.04 189.915 8.09 190.045 ;
		RECT	10.26 189.915 10.31 190.045 ;
		RECT	11.565 189.915 11.615 190.045 ;
		RECT	1.585 189.955 1.715 190.005 ;
		RECT	1.88 189.955 2.01 190.005 ;
		RECT	5.01 189.955 5.14 190.005 ;
		RECT	9.815 189.955 9.945 190.005 ;
		RECT	0.9 190.46 0.95 190.59 ;
		RECT	1.44 190.46 1.49 190.59 ;
		RECT	3.025 190.46 3.075 190.59 ;
		RECT	3.155 190.46 3.205 190.59 ;
		RECT	6.605 190.46 6.655 190.59 ;
		RECT	7.265 190.46 7.315 190.59 ;
		RECT	12.095 190.46 12.145 190.59 ;
		RECT	12.355 190.46 12.405 190.59 ;
		RECT	13.06 190.46 13.11 190.59 ;
		RECT	14.545 190.46 14.595 190.59 ;
		RECT	4.34 190.5 4.47 190.55 ;
		RECT	6.175 190.5 6.305 190.55 ;
		RECT	8.85 190.5 8.98 190.55 ;
		RECT	9.27 190.5 9.4 190.55 ;
		RECT	2.11 190.915 2.16 191.045 ;
		RECT	5.41 190.915 5.46 191.045 ;
		RECT	6.44 190.915 6.49 191.045 ;
		RECT	9.495 190.915 9.545 191.045 ;
		RECT	13.33 190.915 13.38 191.045 ;
		RECT	15.065 190.915 15.115 191.045 ;
		RECT	14.875 190.92 14.925 191.05 ;
		RECT	3.56 190.955 3.69 191.005 ;
		RECT	4.575 191.41 4.625 191.54 ;
		RECT	7.035 191.41 7.085 191.54 ;
		RECT	12.225 191.41 12.275 191.54 ;
		RECT	13.195 191.41 13.245 191.54 ;
		RECT	2.11 191.9 2.16 192.03 ;
		RECT	5.41 191.9 5.46 192.03 ;
		RECT	6.44 191.9 6.49 192.03 ;
		RECT	9.495 191.9 9.545 192.03 ;
		RECT	13.33 191.9 13.38 192.03 ;
		RECT	14.875 191.9 14.925 192.03 ;
		RECT	15.065 191.9 15.115 192.03 ;
		RECT	3.56 191.94 3.69 191.99 ;
		RECT	14.83 192.185 14.96 192.235 ;
		RECT	15.065 192.185 15.115 192.235 ;
		RECT	4.575 192.39 4.625 192.52 ;
		RECT	7.035 192.39 7.085 192.52 ;
		RECT	2.72 192.885 2.77 193.015 ;
		RECT	9.1 192.885 9.15 193.015 ;
		RECT	10.81 192.885 10.86 193.015 ;
		RECT	0.9 193.375 0.95 193.505 ;
		RECT	1.44 193.375 1.49 193.505 ;
		RECT	3.025 193.375 3.075 193.505 ;
		RECT	3.155 193.375 3.205 193.505 ;
		RECT	6.605 193.375 6.655 193.505 ;
		RECT	7.265 193.375 7.315 193.505 ;
		RECT	12.095 193.375 12.145 193.505 ;
		RECT	12.355 193.375 12.405 193.505 ;
		RECT	13.06 193.375 13.11 193.505 ;
		RECT	14.545 193.375 14.595 193.505 ;
		RECT	4.34 193.415 4.47 193.465 ;
		RECT	6.175 193.415 6.305 193.465 ;
		RECT	8.85 193.415 8.98 193.465 ;
		RECT	9.27 193.415 9.4 193.465 ;
		RECT	2.4 193.87 2.45 194 ;
		RECT	2.55 193.87 2.6 194 ;
		RECT	2.86 193.87 2.91 194 ;
		RECT	3.79 193.87 3.84 194 ;
		RECT	4.055 193.87 4.105 194 ;
		RECT	5.575 193.87 5.625 194 ;
		RECT	6.76 193.87 6.81 194 ;
		RECT	8.04 193.87 8.09 194 ;
		RECT	10.26 193.87 10.31 194 ;
		RECT	11.565 193.87 11.615 194 ;
		RECT	1.585 193.91 1.715 193.96 ;
		RECT	1.88 193.91 2.01 193.96 ;
		RECT	5.01 193.91 5.14 193.96 ;
		RECT	0.9 194.36 0.95 194.49 ;
		RECT	1.44 194.36 1.49 194.49 ;
		RECT	3.025 194.36 3.075 194.49 ;
		RECT	3.155 194.36 3.205 194.49 ;
		RECT	6.605 194.36 6.655 194.49 ;
		RECT	7.265 194.36 7.315 194.49 ;
		RECT	12.095 194.36 12.145 194.49 ;
		RECT	12.355 194.36 12.405 194.49 ;
		RECT	13.06 194.36 13.11 194.49 ;
		RECT	14.545 194.36 14.595 194.49 ;
		RECT	4.34 194.4 4.47 194.45 ;
		RECT	6.175 194.4 6.305 194.45 ;
		RECT	8.85 194.4 8.98 194.45 ;
		RECT	9.27 194.4 9.4 194.45 ;
		RECT	2.11 194.855 2.16 194.985 ;
		RECT	5.41 194.855 5.46 194.985 ;
		RECT	6.44 194.855 6.49 194.985 ;
		RECT	9.735 194.855 9.785 194.985 ;
		RECT	10.81 194.855 10.86 194.985 ;
		RECT	13.33 194.855 13.38 194.985 ;
		RECT	14.875 194.855 14.925 194.985 ;
		RECT	15.07 194.855 15.12 194.985 ;
		RECT	3.56 194.895 3.69 194.945 ;
		RECT	4.575 195.345 4.625 195.475 ;
		RECT	2.11 195.835 2.16 195.965 ;
		RECT	5.41 195.835 5.46 195.965 ;
		RECT	6.44 195.835 6.49 195.965 ;
		RECT	9.735 195.835 9.785 195.965 ;
		RECT	10.07 195.835 10.12 195.965 ;
		RECT	10.81 195.835 10.86 195.965 ;
		RECT	13.33 195.835 13.38 195.965 ;
		RECT	14.875 195.835 14.925 195.965 ;
		RECT	15.07 195.835 15.12 195.965 ;
		RECT	3.56 195.875 3.69 195.925 ;
		RECT	0.9 196.33 0.95 196.46 ;
		RECT	1.44 196.33 1.49 196.46 ;
		RECT	3.025 196.33 3.075 196.46 ;
		RECT	3.155 196.33 3.205 196.46 ;
		RECT	6.605 196.33 6.655 196.46 ;
		RECT	7.265 196.33 7.315 196.46 ;
		RECT	12.095 196.33 12.145 196.46 ;
		RECT	12.355 196.33 12.405 196.46 ;
		RECT	13.06 196.33 13.11 196.46 ;
		RECT	14.545 196.33 14.595 196.46 ;
		RECT	4.34 196.37 4.47 196.42 ;
		RECT	6.175 196.37 6.305 196.42 ;
		RECT	8.85 196.37 8.98 196.42 ;
		RECT	9.27 196.37 9.4 196.42 ;
		RECT	2.11 196.82 2.16 196.95 ;
		RECT	5.41 196.82 5.46 196.95 ;
		RECT	6.44 196.82 6.49 196.95 ;
		RECT	10.07 196.82 10.12 196.95 ;
		RECT	10.81 196.82 10.86 196.95 ;
		RECT	13.33 196.82 13.38 196.95 ;
		RECT	14.87 196.82 14.92 196.95 ;
		RECT	15.065 196.82 15.115 196.95 ;
		RECT	3.56 196.86 3.69 196.91 ;
		RECT	0.9 197.31 0.95 197.44 ;
		RECT	1.44 197.31 1.49 197.44 ;
		RECT	3.025 197.31 3.075 197.44 ;
		RECT	3.155 197.31 3.205 197.44 ;
		RECT	6.605 197.31 6.655 197.44 ;
		RECT	7.265 197.31 7.315 197.44 ;
		RECT	12.095 197.31 12.145 197.44 ;
		RECT	12.355 197.31 12.405 197.44 ;
		RECT	13.06 197.31 13.11 197.44 ;
		RECT	14.545 197.31 14.595 197.44 ;
		RECT	4.34 197.35 4.47 197.4 ;
		RECT	6.175 197.35 6.305 197.4 ;
		RECT	8.85 197.35 8.98 197.4 ;
		RECT	9.27 197.35 9.4 197.4 ;
		RECT	2.4 197.805 2.45 197.935 ;
		RECT	2.55 197.805 2.6 197.935 ;
		RECT	2.86 197.805 2.91 197.935 ;
		RECT	3.79 197.805 3.84 197.935 ;
		RECT	4.055 197.805 4.105 197.935 ;
		RECT	5.575 197.805 5.625 197.935 ;
		RECT	6.76 197.805 6.81 197.935 ;
		RECT	8.04 197.805 8.09 197.935 ;
		RECT	10.26 197.805 10.31 197.935 ;
		RECT	11.565 197.805 11.615 197.935 ;
		RECT	1.585 197.845 1.715 197.895 ;
		RECT	1.88 197.845 2.01 197.895 ;
		RECT	5.01 197.845 5.14 197.895 ;
		RECT	0.9 198.295 0.95 198.425 ;
		RECT	1.44 198.295 1.49 198.425 ;
		RECT	3.025 198.295 3.075 198.425 ;
		RECT	3.155 198.295 3.205 198.425 ;
		RECT	6.605 198.295 6.655 198.425 ;
		RECT	7.265 198.295 7.315 198.425 ;
		RECT	12.095 198.295 12.145 198.425 ;
		RECT	12.355 198.295 12.405 198.425 ;
		RECT	13.06 198.295 13.11 198.425 ;
		RECT	14.545 198.295 14.595 198.425 ;
		RECT	4.34 198.335 4.47 198.385 ;
		RECT	6.175 198.335 6.305 198.385 ;
		RECT	8.85 198.335 8.98 198.385 ;
		RECT	9.27 198.335 9.4 198.385 ;
		RECT	2.11 198.79 2.16 198.92 ;
		RECT	5.41 198.79 5.46 198.92 ;
		RECT	6.44 198.79 6.49 198.92 ;
		RECT	6.915 198.79 6.965 198.92 ;
		RECT	10.81 198.79 10.86 198.92 ;
		RECT	13.19 198.79 13.24 198.92 ;
		RECT	13.33 198.79 13.38 198.92 ;
		RECT	14.87 198.79 14.92 198.92 ;
		RECT	15.065 198.79 15.115 198.92 ;
		RECT	3.56 198.83 3.69 198.88 ;
		RECT	4.575 199.28 4.625 199.41 ;
		RECT	7.375 199.565 7.425 199.615 ;
		RECT	3.56 199.745 3.69 199.795 ;
		RECT	2.11 199.77 2.16 199.9 ;
		RECT	5.41 199.77 5.46 199.9 ;
		RECT	6.44 199.77 6.49 199.9 ;
		RECT	6.915 199.77 6.965 199.9 ;
		RECT	7.555 199.77 7.605 199.9 ;
		RECT	10.81 199.77 10.86 199.9 ;
		RECT	13.33 199.77 13.38 199.9 ;
		RECT	14.87 199.77 14.92 199.9 ;
		RECT	15.065 199.77 15.115 199.9 ;
		RECT	3.56 199.875 3.69 199.925 ;
		RECT	4.575 200.265 4.625 200.395 ;
		RECT	2.11 200.755 2.16 200.885 ;
		RECT	5.41 200.755 5.46 200.885 ;
		RECT	6.44 200.755 6.49 200.885 ;
		RECT	6.915 200.755 6.965 200.885 ;
		RECT	7.555 200.755 7.605 200.885 ;
		RECT	10.81 200.755 10.86 200.885 ;
		RECT	13.33 200.755 13.38 200.885 ;
		RECT	14.87 200.755 14.92 200.885 ;
		RECT	15.065 200.755 15.115 200.885 ;
		RECT	3.56 200.795 3.69 200.845 ;
		RECT	0.9 201.25 0.95 201.38 ;
		RECT	1.44 201.25 1.49 201.38 ;
		RECT	3.025 201.25 3.075 201.38 ;
		RECT	3.155 201.25 3.205 201.38 ;
		RECT	6.605 201.25 6.655 201.38 ;
		RECT	7.215 201.25 7.265 201.38 ;
		RECT	12.095 201.25 12.145 201.38 ;
		RECT	12.355 201.25 12.405 201.38 ;
		RECT	13.06 201.25 13.11 201.38 ;
		RECT	14.545 201.25 14.595 201.38 ;
		RECT	4.34 201.29 4.47 201.34 ;
		RECT	6.175 201.29 6.305 201.34 ;
		RECT	8.85 201.29 8.98 201.34 ;
		RECT	9.27 201.29 9.4 201.34 ;
		RECT	9.855 201.535 9.905 201.585 ;
		RECT	9.855 201.535 9.985 201.585 ;
		RECT	1.585 201.715 1.715 201.765 ;
		RECT	1.88 201.715 2.01 201.765 ;
		RECT	5.01 201.715 5.14 201.765 ;
		RECT	2.4 201.74 2.45 201.87 ;
		RECT	2.55 201.74 2.6 201.87 ;
		RECT	2.86 201.74 2.91 201.87 ;
		RECT	3.79 201.74 3.84 201.87 ;
		RECT	4.055 201.74 4.105 201.87 ;
		RECT	5.575 201.74 5.625 201.87 ;
		RECT	6.76 201.74 6.81 201.87 ;
		RECT	8.04 201.74 8.09 201.87 ;
		RECT	10.26 201.74 10.31 201.87 ;
		RECT	11.565 201.74 11.615 201.87 ;
		RECT	1.585 201.845 1.715 201.895 ;
		RECT	1.88 201.845 2.01 201.895 ;
		RECT	5.01 201.845 5.14 201.895 ;
		RECT	0.62 202.235 0.67 202.365 ;
		RECT	1.16 202.235 1.21 202.365 ;
		RECT	4.19 202.235 4.24 202.365 ;
		RECT	7.73 202.235 7.78 202.365 ;
		RECT	14.68 202.235 14.73 202.365 ;
		RECT	2.11 202.73 2.16 202.86 ;
		RECT	5.41 202.73 5.46 202.86 ;
		RECT	6.44 202.73 6.49 202.86 ;
		RECT	6.915 202.73 6.965 202.86 ;
		RECT	7.555 202.73 7.605 202.86 ;
		RECT	10.81 202.73 10.86 202.86 ;
		RECT	13.33 202.73 13.38 202.86 ;
		RECT	14.875 202.73 14.925 202.86 ;
		RECT	15.07 202.73 15.12 202.86 ;
		RECT	3.56 202.77 3.69 202.82 ;
		RECT	4.575 203.215 4.625 203.345 ;
		RECT	12.225 203.215 12.275 203.345 ;
		RECT	14.44 203.215 14.49 203.345 ;
		RECT	2.11 203.71 2.16 203.84 ;
		RECT	5.41 203.71 5.46 203.84 ;
		RECT	6.44 203.71 6.49 203.84 ;
		RECT	6.915 203.71 6.965 203.84 ;
		RECT	7.555 203.71 7.605 203.84 ;
		RECT	10.81 203.71 10.86 203.84 ;
		RECT	13.33 203.71 13.38 203.84 ;
		RECT	14.875 203.71 14.925 203.84 ;
		RECT	15.07 203.71 15.12 203.84 ;
		RECT	3.56 203.75 3.69 203.8 ;
		RECT	14.34 204.185 14.39 204.315 ;
		RECT	15.21 204.185 15.26 204.315 ;
		RECT	14.215 204.81 14.265 204.94 ;
		RECT	1.625 204.865 1.675 204.995 ;
		RECT	1.92 204.865 1.97 204.995 ;
		RECT	2.4 204.865 2.45 204.995 ;
		RECT	2.55 204.865 2.6 204.995 ;
		RECT	2.86 204.865 2.91 204.995 ;
		RECT	3.79 204.865 3.84 204.995 ;
		RECT	4.055 204.865 4.105 204.995 ;
		RECT	5.05 204.865 5.1 204.995 ;
		RECT	5.575 204.865 5.625 204.995 ;
		RECT	6.76 204.865 6.81 204.995 ;
		RECT	8.04 204.865 8.09 204.995 ;
		RECT	10.26 204.865 10.31 204.995 ;
		RECT	11.565 204.865 11.615 204.995 ;
		RECT	4.34 205.16 4.47 205.21 ;
		RECT	6.175 205.16 6.305 205.21 ;
		RECT	8.85 205.16 8.98 205.21 ;
		RECT	9.27 205.16 9.4 205.21 ;
		RECT	0.9 205.185 0.95 205.315 ;
		RECT	1.44 205.185 1.49 205.315 ;
		RECT	3.025 205.185 3.075 205.315 ;
		RECT	3.155 205.185 3.205 205.315 ;
		RECT	6.605 205.185 6.655 205.315 ;
		RECT	7.215 205.185 7.265 205.315 ;
		RECT	12.095 205.185 12.145 205.315 ;
		RECT	12.355 205.185 12.405 205.315 ;
		RECT	13.06 205.185 13.11 205.315 ;
		RECT	14.545 205.185 14.595 205.315 ;
		RECT	4.34 205.29 4.47 205.34 ;
		RECT	6.175 205.29 6.305 205.34 ;
		RECT	8.85 205.29 8.98 205.34 ;
		RECT	9.27 205.29 9.4 205.34 ;
		RECT	14.44 205.47 14.49 205.52 ;
		RECT	1.585 205.65 1.715 205.7 ;
		RECT	1.88 205.65 2.01 205.7 ;
		RECT	5.01 205.65 5.14 205.7 ;
		RECT	2.4 205.675 2.45 205.805 ;
		RECT	2.55 205.675 2.6 205.805 ;
		RECT	2.86 205.675 2.91 205.805 ;
		RECT	3.79 205.675 3.84 205.805 ;
		RECT	4.055 205.675 4.105 205.805 ;
		RECT	5.575 205.675 5.625 205.805 ;
		RECT	6.76 205.675 6.81 205.805 ;
		RECT	8.04 205.675 8.09 205.805 ;
		RECT	10.26 205.675 10.31 205.805 ;
		RECT	11.565 205.675 11.615 205.805 ;
		RECT	1.585 205.78 1.715 205.83 ;
		RECT	1.88 205.78 2.01 205.83 ;
		RECT	5.01 205.78 5.14 205.83 ;
		RECT	14.44 205.965 14.49 206.015 ;
		RECT	0.9 206.17 0.95 206.3 ;
		RECT	1.44 206.17 1.49 206.3 ;
		RECT	3.025 206.17 3.075 206.3 ;
		RECT	3.155 206.17 3.205 206.3 ;
		RECT	6.605 206.17 6.655 206.3 ;
		RECT	7.215 206.17 7.265 206.3 ;
		RECT	10.66 206.17 10.71 206.3 ;
		RECT	12.095 206.17 12.145 206.3 ;
		RECT	12.355 206.17 12.405 206.3 ;
		RECT	13.06 206.17 13.11 206.3 ;
		RECT	14.545 206.17 14.595 206.3 ;
		RECT	4.34 206.21 4.47 206.26 ;
		RECT	6.175 206.21 6.305 206.26 ;
		RECT	8.85 206.21 8.98 206.26 ;
		RECT	9.27 206.21 9.4 206.26 ;
		RECT	2.11 206.66 2.16 206.79 ;
		RECT	5.41 206.66 5.46 206.79 ;
		RECT	6.44 206.66 6.49 206.79 ;
		RECT	6.915 206.66 6.965 206.79 ;
		RECT	7.555 206.66 7.605 206.79 ;
		RECT	9.65 206.66 9.7 206.79 ;
		RECT	10.81 206.66 10.86 206.79 ;
		RECT	13.33 206.66 13.38 206.79 ;
		RECT	14.875 206.66 14.925 206.79 ;
		RECT	15.07 206.66 15.12 206.79 ;
		RECT	3.56 206.7 3.69 206.75 ;
		RECT	4.575 207.15 4.625 207.28 ;
		RECT	14.44 207.15 14.49 207.28 ;
		RECT	7.73 207.44 7.78 207.49 ;
		RECT	13.195 207.44 13.245 207.49 ;
		RECT	4.575 207.645 4.625 207.775 ;
		RECT	14.44 207.645 14.49 207.775 ;
		RECT	2.11 208.135 2.16 208.265 ;
		RECT	5.41 208.135 5.46 208.265 ;
		RECT	6.44 208.135 6.49 208.265 ;
		RECT	6.915 208.135 6.965 208.265 ;
		RECT	7.555 208.135 7.605 208.265 ;
		RECT	9.65 208.135 9.7 208.265 ;
		RECT	10.81 208.135 10.86 208.265 ;
		RECT	13.33 208.135 13.38 208.265 ;
		RECT	14.875 208.135 14.925 208.265 ;
		RECT	15.07 208.135 15.12 208.265 ;
		RECT	3.56 208.175 3.69 208.225 ;
		RECT	0.9 208.63 0.95 208.76 ;
		RECT	1.44 208.63 1.49 208.76 ;
		RECT	3.025 208.63 3.075 208.76 ;
		RECT	3.155 208.63 3.205 208.76 ;
		RECT	6.605 208.63 6.655 208.76 ;
		RECT	7.215 208.63 7.265 208.76 ;
		RECT	10.66 208.63 10.71 208.76 ;
		RECT	12.095 208.63 12.145 208.76 ;
		RECT	12.355 208.63 12.405 208.76 ;
		RECT	13.06 208.63 13.11 208.76 ;
		RECT	14.545 208.63 14.595 208.76 ;
		RECT	4.34 208.67 4.47 208.72 ;
		RECT	4.76 208.67 4.89 208.72 ;
		RECT	6.175 208.67 6.305 208.72 ;
		RECT	8.85 208.67 8.98 208.72 ;
		RECT	9.27 208.67 9.4 208.72 ;
		RECT	14.44 208.915 14.49 208.965 ;
		RECT	5.01 209.095 5.14 209.145 ;
		RECT	2.4 209.12 2.45 209.25 ;
		RECT	2.55 209.12 2.6 209.25 ;
		RECT	2.86 209.12 2.91 209.25 ;
		RECT	3.79 209.12 3.84 209.25 ;
		RECT	4.055 209.12 4.105 209.25 ;
		RECT	5.575 209.12 5.625 209.25 ;
		RECT	6.76 209.12 6.81 209.25 ;
		RECT	8.04 209.12 8.09 209.25 ;
		RECT	10.26 209.12 10.31 209.25 ;
		RECT	11.565 209.12 11.615 209.25 ;
		RECT	1.585 209.16 1.715 209.21 ;
		RECT	1.88 209.16 2.01 209.21 ;
		RECT	5.01 209.225 5.14 209.275 ;
		RECT	14.44 209.405 14.49 209.455 ;
		RECT	4.34 209.585 4.47 209.635 ;
		RECT	6.175 209.585 6.305 209.635 ;
		RECT	8.85 209.585 8.98 209.635 ;
		RECT	9.27 209.585 9.4 209.635 ;
		RECT	0.9 209.61 0.95 209.74 ;
		RECT	1.44 209.61 1.49 209.74 ;
		RECT	3.025 209.61 3.075 209.74 ;
		RECT	3.155 209.61 3.205 209.74 ;
		RECT	6.605 209.61 6.655 209.74 ;
		RECT	7.215 209.61 7.265 209.74 ;
		RECT	12.095 209.61 12.145 209.74 ;
		RECT	12.355 209.61 12.405 209.74 ;
		RECT	13.06 209.61 13.11 209.74 ;
		RECT	14.545 209.61 14.595 209.74 ;
		RECT	4.34 209.715 4.47 209.765 ;
		RECT	6.175 209.715 6.305 209.765 ;
		RECT	8.85 209.715 8.98 209.765 ;
		RECT	9.27 209.715 9.4 209.765 ;
		RECT	14.215 209.925 14.265 210.055 ;
		RECT	1.625 209.93 1.675 210.06 ;
		RECT	1.92 209.93 1.97 210.06 ;
		RECT	2.4 209.93 2.45 210.06 ;
		RECT	2.55 209.93 2.6 210.06 ;
		RECT	2.86 209.93 2.91 210.06 ;
		RECT	3.79 209.93 3.84 210.06 ;
		RECT	4.055 209.93 4.105 210.06 ;
		RECT	5.05 209.93 5.1 210.06 ;
		RECT	5.575 209.93 5.625 210.06 ;
		RECT	6.76 209.93 6.81 210.06 ;
		RECT	8.04 209.93 8.09 210.06 ;
		RECT	10.26 209.93 10.31 210.06 ;
		RECT	11.565 209.93 11.615 210.06 ;
		RECT	14.34 210.61 14.39 210.74 ;
		RECT	15.21 210.61 15.26 210.74 ;
		RECT	2.11 211.085 2.16 211.215 ;
		RECT	5.41 211.085 5.46 211.215 ;
		RECT	6.915 211.085 6.965 211.215 ;
		RECT	7.555 211.085 7.605 211.215 ;
		RECT	10.81 211.085 10.86 211.215 ;
		RECT	13.33 211.085 13.38 211.215 ;
		RECT	14.87 211.085 14.92 211.215 ;
		RECT	15.065 211.085 15.115 211.215 ;
		RECT	3.56 211.125 3.69 211.175 ;
		RECT	4.575 211.58 4.625 211.71 ;
		RECT	13.195 211.58 13.245 211.71 ;
		RECT	14.44 211.58 14.49 211.71 ;
		RECT	2.11 212.075 2.16 212.205 ;
		RECT	5.41 212.075 5.46 212.205 ;
		RECT	6.915 212.075 6.965 212.205 ;
		RECT	7.555 212.075 7.605 212.205 ;
		RECT	10.81 212.075 10.86 212.205 ;
		RECT	13.33 212.075 13.38 212.205 ;
		RECT	14.87 212.075 14.92 212.205 ;
		RECT	15.065 212.075 15.115 212.205 ;
		RECT	3.56 212.115 3.69 212.165 ;
		RECT	0.625 212.565 0.675 212.695 ;
		RECT	1.16 212.565 1.21 212.695 ;
		RECT	4.19 212.565 4.24 212.695 ;
		RECT	7.73 212.565 7.78 212.695 ;
		RECT	14.68 212.565 14.73 212.695 ;
		RECT	7.39 212.85 7.44 212.9 ;
		RECT	1.585 213.03 1.715 213.08 ;
		RECT	1.88 213.03 2.01 213.08 ;
		RECT	5.01 213.03 5.14 213.08 ;
		RECT	2.4 213.055 2.45 213.185 ;
		RECT	2.55 213.055 2.6 213.185 ;
		RECT	2.86 213.055 2.91 213.185 ;
		RECT	3.79 213.055 3.84 213.185 ;
		RECT	4.055 213.055 4.105 213.185 ;
		RECT	5.575 213.055 5.625 213.185 ;
		RECT	6.76 213.055 6.81 213.185 ;
		RECT	8.04 213.055 8.09 213.185 ;
		RECT	10.26 213.055 10.31 213.185 ;
		RECT	11.565 213.055 11.615 213.185 ;
		RECT	1.585 213.16 1.715 213.21 ;
		RECT	1.88 213.16 2.01 213.21 ;
		RECT	5.01 213.16 5.14 213.21 ;
		RECT	0.9 213.55 0.95 213.68 ;
		RECT	1.44 213.55 1.49 213.68 ;
		RECT	3.025 213.55 3.075 213.68 ;
		RECT	3.155 213.55 3.205 213.68 ;
		RECT	6.605 213.55 6.655 213.68 ;
		RECT	7.215 213.55 7.265 213.68 ;
		RECT	12.095 213.55 12.145 213.68 ;
		RECT	12.355 213.55 12.405 213.68 ;
		RECT	13.06 213.55 13.11 213.68 ;
		RECT	14.545 213.55 14.595 213.68 ;
		RECT	4.34 213.59 4.47 213.64 ;
		RECT	6.175 213.59 6.305 213.64 ;
		RECT	8.85 213.59 8.98 213.64 ;
		RECT	9.27 213.59 9.4 213.64 ;
		RECT	2.11 214.04 2.16 214.17 ;
		RECT	5.41 214.04 5.46 214.17 ;
		RECT	6.915 214.04 6.965 214.17 ;
		RECT	7.555 214.04 7.605 214.17 ;
		RECT	10.81 214.04 10.86 214.17 ;
		RECT	13.33 214.04 13.38 214.17 ;
		RECT	14.87 214.04 14.92 214.17 ;
		RECT	15.065 214.04 15.115 214.17 ;
		RECT	3.56 214.08 3.69 214.13 ;
		RECT	4.575 214.535 4.625 214.665 ;
		RECT	13.195 214.535 13.245 214.665 ;
		RECT	14.44 214.535 14.49 214.665 ;
		RECT	3.56 215 3.69 215.05 ;
		RECT	2.11 215.025 2.16 215.155 ;
		RECT	5.41 215.025 5.46 215.155 ;
		RECT	6.915 215.025 6.965 215.155 ;
		RECT	7.555 215.025 7.605 215.155 ;
		RECT	10.81 215.025 10.86 215.155 ;
		RECT	13.33 215.025 13.38 215.155 ;
		RECT	14.87 215.025 14.92 215.155 ;
		RECT	15.065 215.025 15.115 215.155 ;
		RECT	3.56 215.13 3.69 215.18 ;
		RECT	7.39 215.31 7.44 215.36 ;
		RECT	4.575 215.515 4.625 215.645 ;
		RECT	13.195 215.515 13.245 215.645 ;
		RECT	2.11 216.01 2.16 216.14 ;
		RECT	5.41 216.01 5.46 216.14 ;
		RECT	6.915 216.01 6.965 216.14 ;
		RECT	10.81 216.01 10.86 216.14 ;
		RECT	13.33 216.01 13.38 216.14 ;
		RECT	14.87 216.01 14.92 216.14 ;
		RECT	15.065 216.01 15.115 216.14 ;
		RECT	3.56 216.05 3.69 216.1 ;
		RECT	0.9 216.5 0.95 216.63 ;
		RECT	1.44 216.5 1.49 216.63 ;
		RECT	3.025 216.5 3.075 216.63 ;
		RECT	3.155 216.5 3.205 216.63 ;
		RECT	6.605 216.5 6.655 216.63 ;
		RECT	7.265 216.5 7.315 216.63 ;
		RECT	12.095 216.5 12.145 216.63 ;
		RECT	12.355 216.5 12.405 216.63 ;
		RECT	13.06 216.5 13.11 216.63 ;
		RECT	14.545 216.5 14.595 216.63 ;
		RECT	4.34 216.54 4.47 216.59 ;
		RECT	6.175 216.54 6.305 216.59 ;
		RECT	8.85 216.54 8.98 216.59 ;
		RECT	9.27 216.54 9.4 216.59 ;
		RECT	2.4 216.995 2.45 217.125 ;
		RECT	2.55 216.995 2.6 217.125 ;
		RECT	2.86 216.995 2.91 217.125 ;
		RECT	3.79 216.995 3.84 217.125 ;
		RECT	4.055 216.995 4.105 217.125 ;
		RECT	6.76 216.995 6.81 217.125 ;
		RECT	8.04 216.995 8.09 217.125 ;
		RECT	10.26 216.995 10.31 217.125 ;
		RECT	11.565 216.995 11.615 217.125 ;
		RECT	1.585 217.035 1.715 217.085 ;
		RECT	1.88 217.035 2.01 217.085 ;
		RECT	5.01 217.035 5.14 217.085 ;
		RECT	9.79 217.035 9.92 217.085 ;
		RECT	0.9 217.485 0.95 217.615 ;
		RECT	1.44 217.485 1.49 217.615 ;
		RECT	3.025 217.485 3.075 217.615 ;
		RECT	3.155 217.485 3.205 217.615 ;
		RECT	6.605 217.485 6.655 217.615 ;
		RECT	7.265 217.485 7.315 217.615 ;
		RECT	12.095 217.485 12.145 217.615 ;
		RECT	12.355 217.485 12.405 217.615 ;
		RECT	13.06 217.485 13.11 217.615 ;
		RECT	14.545 217.485 14.595 217.615 ;
		RECT	4.34 217.525 4.47 217.575 ;
		RECT	6.175 217.525 6.305 217.575 ;
		RECT	8.85 217.525 8.98 217.575 ;
		RECT	9.27 217.525 9.4 217.575 ;
		RECT	2.11 217.975 2.16 218.105 ;
		RECT	5.41 217.975 5.46 218.105 ;
		RECT	6.915 217.975 6.965 218.105 ;
		RECT	10.81 217.975 10.86 218.105 ;
		RECT	13.33 217.975 13.38 218.105 ;
		RECT	14.87 217.975 14.92 218.105 ;
		RECT	15.065 217.975 15.115 218.105 ;
		RECT	3.56 218.015 3.69 218.065 ;
		RECT	0.9 218.47 0.95 218.6 ;
		RECT	1.44 218.47 1.49 218.6 ;
		RECT	3.025 218.47 3.075 218.6 ;
		RECT	3.155 218.47 3.205 218.6 ;
		RECT	6.605 218.47 6.655 218.6 ;
		RECT	7.265 218.47 7.315 218.6 ;
		RECT	12.095 218.47 12.145 218.6 ;
		RECT	12.355 218.47 12.405 218.6 ;
		RECT	13.06 218.47 13.11 218.6 ;
		RECT	14.545 218.47 14.595 218.6 ;
		RECT	4.34 218.51 4.47 218.56 ;
		RECT	6.175 218.51 6.305 218.56 ;
		RECT	8.85 218.51 8.98 218.56 ;
		RECT	9.27 218.51 9.4 218.56 ;
		RECT	2.11 218.96 2.16 219.09 ;
		RECT	5.41 218.96 5.46 219.09 ;
		RECT	6.915 218.96 6.965 219.09 ;
		RECT	10.81 218.96 10.86 219.09 ;
		RECT	13.33 218.96 13.38 219.09 ;
		RECT	14.87 218.96 14.92 219.09 ;
		RECT	15.065 218.96 15.115 219.09 ;
		RECT	3.56 219 3.69 219.05 ;
		RECT	13.195 219.445 13.245 219.575 ;
		RECT	4.575 219.455 4.625 219.585 ;
		RECT	2.11 219.945 2.16 220.075 ;
		RECT	5.41 219.945 5.46 220.075 ;
		RECT	6.915 219.945 6.965 220.075 ;
		RECT	10.81 219.945 10.86 220.075 ;
		RECT	13.33 219.945 13.38 220.075 ;
		RECT	14.87 219.945 14.92 220.075 ;
		RECT	15.065 219.945 15.115 220.075 ;
		RECT	3.56 219.985 3.69 220.035 ;
		RECT	0.9 220.435 0.95 220.565 ;
		RECT	1.44 220.435 1.49 220.565 ;
		RECT	3.025 220.435 3.075 220.565 ;
		RECT	3.155 220.435 3.205 220.565 ;
		RECT	6.605 220.435 6.655 220.565 ;
		RECT	7.265 220.435 7.315 220.565 ;
		RECT	12.095 220.435 12.145 220.565 ;
		RECT	12.355 220.435 12.405 220.565 ;
		RECT	13.06 220.435 13.11 220.565 ;
		RECT	14.545 220.435 14.595 220.565 ;
		RECT	4.34 220.475 4.47 220.525 ;
		RECT	6.175 220.475 6.305 220.525 ;
		RECT	8.85 220.475 8.98 220.525 ;
		RECT	9.27 220.475 9.4 220.525 ;
		RECT	14.83 220.72 14.96 220.77 ;
		RECT	15.065 220.72 15.115 220.77 ;
		RECT	1.585 220.905 1.715 220.955 ;
		RECT	1.88 220.905 2.01 220.955 ;
		RECT	5.01 220.905 5.14 220.955 ;
		RECT	9.815 220.905 9.945 220.955 ;
		RECT	2.4 220.93 2.45 221.06 ;
		RECT	2.55 220.93 2.6 221.06 ;
		RECT	2.86 220.93 2.91 221.06 ;
		RECT	3.79 220.93 3.84 221.06 ;
		RECT	4.055 220.93 4.105 221.06 ;
		RECT	6.76 220.93 6.81 221.06 ;
		RECT	8.04 220.93 8.09 221.06 ;
		RECT	10.26 220.93 10.31 221.06 ;
		RECT	11.565 220.93 11.615 221.06 ;
		RECT	1.585 221.035 1.715 221.085 ;
		RECT	1.88 221.035 2.01 221.085 ;
		RECT	5.01 221.035 5.14 221.085 ;
		RECT	9.815 221.035 9.945 221.085 ;
		RECT	0.905 221.215 1.035 221.265 ;
		RECT	1.355 221.215 1.485 221.265 ;
		RECT	3.05 221.215 3.18 221.265 ;
		RECT	0.9 221.42 0.95 221.55 ;
		RECT	1.44 221.42 1.49 221.55 ;
		RECT	3.025 221.42 3.075 221.55 ;
		RECT	3.155 221.42 3.205 221.55 ;
		RECT	6.605 221.42 6.655 221.55 ;
		RECT	7.265 221.42 7.315 221.55 ;
		RECT	12.095 221.42 12.145 221.55 ;
		RECT	12.355 221.42 12.405 221.55 ;
		RECT	13.06 221.42 13.11 221.55 ;
		RECT	14.545 221.42 14.595 221.55 ;
		RECT	4.34 221.46 4.47 221.51 ;
		RECT	6.175 221.46 6.305 221.51 ;
		RECT	8.85 221.46 8.98 221.51 ;
		RECT	9.27 221.46 9.4 221.51 ;
		RECT	2.72 221.915 2.77 222.045 ;
		RECT	9.1 221.915 9.15 222.045 ;
		RECT	10.81 221.915 10.86 222.045 ;
		RECT	4.575 222.405 4.625 222.535 ;
		RECT	3.56 222.87 3.69 222.92 ;
		RECT	2.11 222.895 2.16 223.025 ;
		RECT	5.41 222.895 5.46 223.025 ;
		RECT	6.915 222.895 6.965 223.025 ;
		RECT	12.23 222.895 12.28 223.025 ;
		RECT	13.33 222.895 13.38 223.025 ;
		RECT	14.87 222.895 14.92 223.025 ;
		RECT	15.065 222.895 15.115 223.025 ;
		RECT	3.56 223 3.69 223.05 ;
		RECT	4.575 223.355 4.625 223.485 ;
		RECT	13.195 223.355 13.245 223.485 ;
		RECT	2.11 223.88 2.16 224.01 ;
		RECT	5.41 223.88 5.46 224.01 ;
		RECT	6.915 223.88 6.965 224.01 ;
		RECT	12.23 223.88 12.28 224.01 ;
		RECT	13.33 223.88 13.38 224.01 ;
		RECT	14.87 223.88 14.92 224.01 ;
		RECT	15.065 223.88 15.115 224.01 ;
		RECT	3.56 223.92 3.69 223.97 ;
		RECT	0.9 224.34 0.95 224.47 ;
		RECT	1.44 224.34 1.49 224.47 ;
		RECT	3.025 224.34 3.075 224.47 ;
		RECT	3.155 224.34 3.205 224.47 ;
		RECT	6.605 224.34 6.655 224.47 ;
		RECT	7.265 224.34 7.315 224.47 ;
		RECT	12.095 224.34 12.145 224.47 ;
		RECT	12.355 224.34 12.405 224.47 ;
		RECT	13.06 224.34 13.11 224.47 ;
		RECT	14.545 224.34 14.595 224.47 ;
		RECT	4.34 224.38 4.47 224.43 ;
		RECT	6.175 224.38 6.305 224.43 ;
		RECT	8.85 224.38 8.98 224.43 ;
		RECT	9.27 224.38 9.4 224.43 ;
		RECT	2.4 224.88 2.45 225.01 ;
		RECT	2.55 224.88 2.6 225.01 ;
		RECT	3.79 224.88 3.84 225.01 ;
		RECT	4.055 224.88 4.105 225.01 ;
		RECT	6.76 224.88 6.81 225.01 ;
		RECT	8.04 224.88 8.09 225.01 ;
		RECT	10.26 224.88 10.31 225.01 ;
		RECT	11.565 224.88 11.615 225.01 ;
		RECT	1.585 224.92 1.715 224.97 ;
		RECT	1.88 224.92 2.01 224.97 ;
		RECT	5.01 224.92 5.14 224.97 ;
		RECT	9.815 224.92 9.945 224.97 ;
		RECT	13.195 225.155 13.245 225.205 ;
		RECT	1.585 225.33 1.715 225.38 ;
		RECT	1.88 225.33 2.01 225.38 ;
		RECT	5.01 225.33 5.14 225.38 ;
		RECT	9.815 225.33 9.945 225.38 ;
		RECT	2.4 225.355 2.45 225.485 ;
		RECT	2.55 225.355 2.6 225.485 ;
		RECT	3.79 225.355 3.84 225.485 ;
		RECT	4.055 225.355 4.105 225.485 ;
		RECT	6.76 225.355 6.81 225.485 ;
		RECT	8.04 225.355 8.09 225.485 ;
		RECT	10.26 225.355 10.31 225.485 ;
		RECT	11.565 225.355 11.615 225.485 ;
		RECT	14.215 225.355 14.265 225.485 ;
		RECT	1.585 225.46 1.715 225.51 ;
		RECT	1.88 225.46 2.01 225.51 ;
		RECT	5.01 225.46 5.14 225.51 ;
		RECT	9.815 225.46 9.945 225.51 ;
		RECT	2.11 225.85 2.16 225.98 ;
		RECT	5.41 225.85 5.46 225.98 ;
		RECT	6.915 225.85 6.965 225.98 ;
		RECT	9.515 225.85 9.565 225.98 ;
		RECT	12.23 225.85 12.28 225.98 ;
		RECT	13.33 225.85 13.38 225.98 ;
		RECT	14.87 225.85 14.92 225.98 ;
		RECT	15.065 225.85 15.115 225.98 ;
		RECT	3.56 225.89 3.69 225.94 ;
		RECT	13.195 226.135 13.245 226.185 ;
		RECT	0.9 226.34 0.95 226.47 ;
		RECT	1.44 226.34 1.49 226.47 ;
		RECT	3.025 226.34 3.075 226.47 ;
		RECT	3.155 226.34 3.205 226.47 ;
		RECT	6.605 226.34 6.655 226.47 ;
		RECT	7.265 226.34 7.315 226.47 ;
		RECT	12.095 226.34 12.145 226.47 ;
		RECT	12.355 226.34 12.405 226.47 ;
		RECT	13.06 226.34 13.11 226.47 ;
		RECT	14.545 226.34 14.595 226.47 ;
		RECT	4.34 226.38 4.47 226.43 ;
		RECT	6.175 226.38 6.305 226.43 ;
		RECT	8.85 226.38 8.98 226.43 ;
		RECT	9.27 226.38 9.4 226.43 ;
		RECT	2.11 226.835 2.16 226.965 ;
		RECT	5.41 226.835 5.46 226.965 ;
		RECT	6.915 226.835 6.965 226.965 ;
		RECT	9.515 226.835 9.565 226.965 ;
		RECT	12.23 226.835 12.28 226.965 ;
		RECT	13.33 226.835 13.38 226.965 ;
		RECT	14.87 226.835 14.92 226.965 ;
		RECT	15.065 226.835 15.115 226.965 ;
		RECT	3.56 226.875 3.69 226.925 ;
		RECT	1.585 227.12 1.715 227.17 ;
		RECT	1.88 227.12 2.01 227.17 ;
		RECT	5.01 227.12 5.14 227.17 ;
		RECT	9.815 227.12 9.945 227.17 ;
		RECT	2.4 227.145 2.45 227.275 ;
		RECT	2.55 227.145 2.6 227.275 ;
		RECT	3.79 227.145 3.84 227.275 ;
		RECT	4.055 227.145 4.105 227.275 ;
		RECT	6.76 227.145 6.81 227.275 ;
		RECT	8.04 227.145 8.09 227.275 ;
		RECT	10.26 227.145 10.31 227.275 ;
		RECT	11.565 227.145 11.615 227.275 ;
		RECT	1.585 227.25 1.715 227.3 ;
		RECT	1.88 227.25 2.01 227.3 ;
		RECT	5.01 227.25 5.14 227.3 ;
		RECT	9.815 227.25 9.945 227.3 ;
		RECT	14.34 227.625 14.39 227.755 ;
		RECT	2.72 227.855 2.77 227.985 ;
		RECT	9.1 227.855 9.15 227.985 ;
		RECT	10.81 227.855 10.86 227.985 ;
		RECT	0.62 228.085 0.67 228.215 ;
		RECT	1.16 228.085 1.21 228.215 ;
		RECT	4.19 228.085 4.24 228.215 ;
		RECT	7.73 228.085 7.78 228.215 ;
		RECT	14.68 228.085 14.73 228.215 ;
		RECT	1.625 228.315 1.675 228.445 ;
		RECT	1.92 228.315 1.97 228.445 ;
		RECT	2.4 228.315 2.45 228.445 ;
		RECT	2.55 228.315 2.6 228.445 ;
		RECT	3.79 228.315 3.84 228.445 ;
		RECT	4.055 228.315 4.105 228.445 ;
		RECT	5.05 228.315 5.1 228.445 ;
		RECT	6.76 228.315 6.81 228.445 ;
		RECT	8.04 228.315 8.09 228.445 ;
		RECT	9.855 228.315 9.905 228.445 ;
		RECT	10.26 228.315 10.31 228.445 ;
		RECT	11.565 228.315 11.615 228.445 ;
		RECT	0.435 187.965 0.485 188.095 ;
		RECT	0.435 188.945 0.485 189.075 ;
		RECT	0.435 190.915 0.485 191.045 ;
		RECT	0.435 191.9 0.485 192.03 ;
		RECT	0.435 194.855 0.485 194.985 ;
		RECT	0.435 195.835 0.485 195.965 ;
		RECT	0.435 196.82 0.485 196.95 ;
		RECT	0.435 198.79 0.485 198.92 ;
		RECT	0.17 199.57 0.22 199.62 ;
		RECT	0.435 199.77 0.485 199.9 ;
		RECT	0.435 200.755 0.485 200.885 ;
		RECT	0.18 201.535 0.23 201.585 ;
		RECT	0.435 202.73 0.485 202.86 ;
		RECT	0.435 203.71 0.485 203.84 ;
		RECT	0.435 206.66 0.485 206.79 ;
		RECT	0.435 208.135 0.485 208.265 ;
		RECT	0.435 211.085 0.485 211.215 ;
		RECT	0.435 212.075 0.485 212.205 ;
		RECT	0.18 212.85 0.23 212.9 ;
		RECT	0.435 214.04 0.485 214.17 ;
		RECT	0.435 215.025 0.485 215.155 ;
		RECT	0.17 215.31 0.22 215.36 ;
		RECT	0.435 216.01 0.485 216.14 ;
		RECT	0.435 217.975 0.485 218.105 ;
		RECT	0.435 218.96 0.485 219.09 ;
		RECT	0.435 219.945 0.485 220.075 ;
		RECT	0.17 221.215 0.22 221.265 ;
		RECT	0.435 222.2 0.485 222.25 ;
		RECT	0.435 222.69 0.485 222.74 ;
		RECT	0.435 222.895 0.485 223.025 ;
		RECT	0.435 223.88 0.485 224.01 ;
		RECT	0.435 225.85 0.485 225.98 ;
		RECT	0.435 226.835 0.485 226.965 ;
		RECT	2.11 186.415 2.16 186.545 ;
		RECT	3.6 186.415 3.65 186.545 ;
		RECT	5.41 186.415 5.46 186.545 ;
		RECT	13.33 186.415 13.38 186.545 ;
		RECT	2.11 187.58 2.16 187.71 ;
		RECT	5.41 187.58 5.46 187.71 ;
		RECT	9.495 187.58 9.545 187.71 ;
		RECT	13.33 187.58 13.38 187.71 ;
		RECT	2.4 187.965 2.45 188.095 ;
		RECT	2.55 187.965 2.6 188.095 ;
		RECT	3.79 187.965 3.84 188.095 ;
		RECT	4.055 187.965 4.105 188.095 ;
		RECT	5.575 187.965 5.625 188.095 ;
		RECT	6.76 187.965 6.81 188.095 ;
		RECT	8.04 187.965 8.09 188.095 ;
		RECT	10.26 187.965 10.31 188.095 ;
		RECT	11.565 187.965 11.615 188.095 ;
		RECT	2.4 188.945 2.45 189.075 ;
		RECT	2.55 188.945 2.6 189.075 ;
		RECT	3.79 188.945 3.84 189.075 ;
		RECT	4.055 188.945 4.105 189.075 ;
		RECT	5.575 188.945 5.625 189.075 ;
		RECT	6.76 188.945 6.81 189.075 ;
		RECT	8.04 188.945 8.09 189.075 ;
		RECT	10.26 188.945 10.31 189.075 ;
		RECT	11.565 188.945 11.615 189.075 ;
		RECT	2.11 189.445 2.16 189.575 ;
		RECT	3.56 189.42 3.69 189.6 ;
		RECT	5.41 189.445 5.46 189.575 ;
		RECT	6.44 189.445 6.49 189.575 ;
		RECT	9.495 189.445 9.545 189.575 ;
		RECT	2.11 189.915 2.16 190.045 ;
		RECT	3.56 189.89 3.69 190.07 ;
		RECT	5.41 189.915 5.46 190.045 ;
		RECT	6.44 189.915 6.49 190.045 ;
		RECT	9.495 189.915 9.545 190.045 ;
		RECT	13.33 189.915 13.38 190.045 ;
		RECT	2.4 190.915 2.45 191.045 ;
		RECT	2.55 190.915 2.6 191.045 ;
		RECT	3.79 190.915 3.84 191.045 ;
		RECT	4.055 190.915 4.105 191.045 ;
		RECT	5.575 190.915 5.625 191.045 ;
		RECT	6.76 190.915 6.81 191.045 ;
		RECT	8.04 190.915 8.09 191.045 ;
		RECT	10.26 190.915 10.31 191.045 ;
		RECT	11.565 190.915 11.615 191.045 ;
		RECT	2.4 191.9 2.45 192.03 ;
		RECT	2.55 191.9 2.6 192.03 ;
		RECT	3.79 191.9 3.84 192.03 ;
		RECT	4.055 191.9 4.105 192.03 ;
		RECT	5.575 191.9 5.625 192.03 ;
		RECT	6.76 191.9 6.81 192.03 ;
		RECT	8.04 191.9 8.09 192.03 ;
		RECT	10.26 191.9 10.31 192.03 ;
		RECT	11.565 191.9 11.615 192.03 ;
		RECT	2.11 193.87 2.16 194 ;
		RECT	5.41 193.87 5.46 194 ;
		RECT	6.44 193.87 6.49 194 ;
		RECT	13.33 193.87 13.38 194 ;
		RECT	2.4 194.855 2.45 194.985 ;
		RECT	2.55 194.855 2.6 194.985 ;
		RECT	2.86 194.855 2.91 194.985 ;
		RECT	3.79 194.855 3.84 194.985 ;
		RECT	4.055 194.855 4.105 194.985 ;
		RECT	5.575 194.855 5.625 194.985 ;
		RECT	6.76 194.855 6.81 194.985 ;
		RECT	8.04 194.855 8.09 194.985 ;
		RECT	10.26 194.855 10.31 194.985 ;
		RECT	11.565 194.855 11.615 194.985 ;
		RECT	2.4 195.835 2.45 195.965 ;
		RECT	2.55 195.835 2.6 195.965 ;
		RECT	2.86 195.835 2.91 195.965 ;
		RECT	3.79 195.835 3.84 195.965 ;
		RECT	4.055 195.835 4.105 195.965 ;
		RECT	5.575 195.835 5.625 195.965 ;
		RECT	6.76 195.835 6.81 195.965 ;
		RECT	8.04 195.835 8.09 195.965 ;
		RECT	10.26 195.835 10.31 195.965 ;
		RECT	11.565 195.835 11.615 195.965 ;
		RECT	2.4 196.82 2.45 196.95 ;
		RECT	2.55 196.82 2.6 196.95 ;
		RECT	2.86 196.82 2.91 196.95 ;
		RECT	3.79 196.82 3.84 196.95 ;
		RECT	4.055 196.82 4.105 196.95 ;
		RECT	5.575 196.82 5.625 196.95 ;
		RECT	6.76 196.82 6.81 196.95 ;
		RECT	8.04 196.82 8.09 196.95 ;
		RECT	10.26 196.82 10.31 196.95 ;
		RECT	11.565 196.82 11.615 196.95 ;
		RECT	2.11 197.805 2.16 197.935 ;
		RECT	5.41 197.805 5.46 197.935 ;
		RECT	6.44 197.805 6.49 197.935 ;
		RECT	10.07 197.805 10.12 197.935 ;
		RECT	10.81 197.805 10.86 197.935 ;
		RECT	13.33 197.805 13.38 197.935 ;
		RECT	2.4 198.79 2.45 198.92 ;
		RECT	2.55 198.79 2.6 198.92 ;
		RECT	2.86 198.79 2.91 198.92 ;
		RECT	3.79 198.79 3.84 198.92 ;
		RECT	4.055 198.79 4.105 198.92 ;
		RECT	5.575 198.79 5.625 198.92 ;
		RECT	6.76 198.79 6.81 198.92 ;
		RECT	8.04 198.79 8.09 198.92 ;
		RECT	10.26 198.79 10.31 198.92 ;
		RECT	11.565 198.79 11.615 198.92 ;
		RECT	2.4 199.77 2.45 199.9 ;
		RECT	2.55 199.77 2.6 199.9 ;
		RECT	2.86 199.77 2.91 199.9 ;
		RECT	3.79 199.77 3.84 199.9 ;
		RECT	4.055 199.77 4.105 199.9 ;
		RECT	5.01 199.745 5.14 199.925 ;
		RECT	5.575 199.77 5.625 199.9 ;
		RECT	6.76 199.77 6.81 199.9 ;
		RECT	8.04 199.77 8.09 199.9 ;
		RECT	10.26 199.77 10.31 199.9 ;
		RECT	11.565 199.77 11.615 199.9 ;
		RECT	2.4 200.755 2.45 200.885 ;
		RECT	2.55 200.755 2.6 200.885 ;
		RECT	2.86 200.755 2.91 200.885 ;
		RECT	3.79 200.755 3.84 200.885 ;
		RECT	4.055 200.755 4.105 200.885 ;
		RECT	5.575 200.755 5.625 200.885 ;
		RECT	6.76 200.755 6.81 200.885 ;
		RECT	8.04 200.755 8.09 200.885 ;
		RECT	10.26 200.755 10.31 200.885 ;
		RECT	11.565 200.755 11.615 200.885 ;
		RECT	2.11 201.74 2.16 201.87 ;
		RECT	3.56 201.715 3.69 201.895 ;
		RECT	5.41 201.74 5.46 201.87 ;
		RECT	6.44 201.74 6.49 201.87 ;
		RECT	6.915 201.74 6.965 201.87 ;
		RECT	7.555 201.74 7.605 201.87 ;
		RECT	10.81 201.74 10.86 201.87 ;
		RECT	13.33 201.74 13.38 201.87 ;
		RECT	14.83 201.715 14.96 201.895 ;
		RECT	2.4 202.73 2.45 202.86 ;
		RECT	2.55 202.73 2.6 202.86 ;
		RECT	2.86 202.73 2.91 202.86 ;
		RECT	3.79 202.73 3.84 202.86 ;
		RECT	4.055 202.73 4.105 202.86 ;
		RECT	5.575 202.73 5.625 202.86 ;
		RECT	6.76 202.73 6.81 202.86 ;
		RECT	8.04 202.73 8.09 202.86 ;
		RECT	10.26 202.73 10.31 202.86 ;
		RECT	11.565 202.73 11.615 202.86 ;
		RECT	2.4 203.71 2.45 203.84 ;
		RECT	2.55 203.71 2.6 203.84 ;
		RECT	2.86 203.71 2.91 203.84 ;
		RECT	3.79 203.71 3.84 203.84 ;
		RECT	4.055 203.71 4.105 203.84 ;
		RECT	5.575 203.71 5.625 203.84 ;
		RECT	6.76 203.71 6.81 203.84 ;
		RECT	8.04 203.71 8.09 203.84 ;
		RECT	10.26 203.71 10.31 203.84 ;
		RECT	11.565 203.71 11.615 203.84 ;
		RECT	2.11 204.865 2.16 204.995 ;
		RECT	3.6 204.865 3.65 204.995 ;
		RECT	5.41 204.865 5.46 204.995 ;
		RECT	6.44 204.865 6.49 204.995 ;
		RECT	6.915 204.865 6.965 204.995 ;
		RECT	7.555 204.865 7.605 204.995 ;
		RECT	9.65 204.865 9.7 204.995 ;
		RECT	10.81 204.865 10.86 204.995 ;
		RECT	2.11 205.675 2.16 205.805 ;
		RECT	3.56 205.65 3.69 205.83 ;
		RECT	5.41 205.675 5.46 205.805 ;
		RECT	6.44 205.675 6.49 205.805 ;
		RECT	6.915 205.675 6.965 205.805 ;
		RECT	7.555 205.675 7.605 205.805 ;
		RECT	9.65 205.675 9.7 205.805 ;
		RECT	10.81 205.675 10.86 205.805 ;
		RECT	13.33 205.675 13.38 205.805 ;
		RECT	2.4 206.66 2.45 206.79 ;
		RECT	2.55 206.66 2.6 206.79 ;
		RECT	2.86 206.66 2.91 206.79 ;
		RECT	3.79 206.66 3.84 206.79 ;
		RECT	4.055 206.66 4.105 206.79 ;
		RECT	5.575 206.66 5.625 206.79 ;
		RECT	6.76 206.66 6.81 206.79 ;
		RECT	8.04 206.66 8.09 206.79 ;
		RECT	10.26 206.66 10.31 206.79 ;
		RECT	11.565 206.66 11.615 206.79 ;
		RECT	2.4 208.135 2.45 208.265 ;
		RECT	2.55 208.135 2.6 208.265 ;
		RECT	2.86 208.135 2.91 208.265 ;
		RECT	3.79 208.135 3.84 208.265 ;
		RECT	4.055 208.135 4.105 208.265 ;
		RECT	5.575 208.135 5.625 208.265 ;
		RECT	6.76 208.135 6.81 208.265 ;
		RECT	8.04 208.135 8.09 208.265 ;
		RECT	10.26 208.135 10.31 208.265 ;
		RECT	11.565 208.135 11.615 208.265 ;
		RECT	2.11 209.12 2.16 209.25 ;
		RECT	3.56 209.095 3.69 209.275 ;
		RECT	5.41 209.12 5.46 209.25 ;
		RECT	6.915 209.12 6.965 209.25 ;
		RECT	7.555 209.12 7.605 209.25 ;
		RECT	9.65 209.12 9.7 209.25 ;
		RECT	10.81 209.12 10.86 209.25 ;
		RECT	13.33 209.12 13.38 209.25 ;
		RECT	2.11 209.93 2.16 210.06 ;
		RECT	3.6 209.93 3.65 210.06 ;
		RECT	5.41 209.93 5.46 210.06 ;
		RECT	6.915 209.93 6.965 210.06 ;
		RECT	7.555 209.93 7.605 210.06 ;
		RECT	9.65 209.93 9.7 210.06 ;
		RECT	10.81 209.93 10.86 210.06 ;
		RECT	2.4 211.085 2.45 211.215 ;
		RECT	2.55 211.085 2.6 211.215 ;
		RECT	2.86 211.085 2.91 211.215 ;
		RECT	3.79 211.085 3.84 211.215 ;
		RECT	4.055 211.085 4.105 211.215 ;
		RECT	5.575 211.085 5.625 211.215 ;
		RECT	6.76 211.085 6.81 211.215 ;
		RECT	8.04 211.085 8.09 211.215 ;
		RECT	10.26 211.085 10.31 211.215 ;
		RECT	11.565 211.085 11.615 211.215 ;
		RECT	2.4 212.075 2.45 212.205 ;
		RECT	2.55 212.075 2.6 212.205 ;
		RECT	2.86 212.075 2.91 212.205 ;
		RECT	3.79 212.075 3.84 212.205 ;
		RECT	4.055 212.075 4.105 212.205 ;
		RECT	5.575 212.075 5.625 212.205 ;
		RECT	6.76 212.075 6.81 212.205 ;
		RECT	8.04 212.075 8.09 212.205 ;
		RECT	10.26 212.075 10.31 212.205 ;
		RECT	11.565 212.075 11.615 212.205 ;
		RECT	2.11 213.055 2.16 213.185 ;
		RECT	3.56 213.03 3.69 213.21 ;
		RECT	5.41 213.055 5.46 213.185 ;
		RECT	6.915 213.055 6.965 213.185 ;
		RECT	7.555 213.055 7.605 213.185 ;
		RECT	10.81 213.055 10.86 213.185 ;
		RECT	13.33 213.055 13.38 213.185 ;
		RECT	14.83 213.03 14.96 213.21 ;
		RECT	2.4 214.04 2.45 214.17 ;
		RECT	2.55 214.04 2.6 214.17 ;
		RECT	2.86 214.04 2.91 214.17 ;
		RECT	3.79 214.04 3.84 214.17 ;
		RECT	4.055 214.04 4.105 214.17 ;
		RECT	5.575 214.04 5.625 214.17 ;
		RECT	6.76 214.04 6.81 214.17 ;
		RECT	8.04 214.04 8.09 214.17 ;
		RECT	10.26 214.04 10.31 214.17 ;
		RECT	11.565 214.04 11.615 214.17 ;
		RECT	2.4 215.025 2.45 215.155 ;
		RECT	2.55 215.025 2.6 215.155 ;
		RECT	2.86 215.025 2.91 215.155 ;
		RECT	3.79 215.025 3.84 215.155 ;
		RECT	4.055 215.025 4.105 215.155 ;
		RECT	5.01 215 5.14 215.18 ;
		RECT	5.575 215.025 5.625 215.155 ;
		RECT	6.76 215.025 6.81 215.155 ;
		RECT	8.04 215.025 8.09 215.155 ;
		RECT	9.79 215 9.92 215.18 ;
		RECT	10.26 215.025 10.31 215.155 ;
		RECT	11.565 215.025 11.615 215.155 ;
		RECT	2.4 216.01 2.45 216.14 ;
		RECT	2.55 216.01 2.6 216.14 ;
		RECT	2.86 216.01 2.91 216.14 ;
		RECT	3.79 216.01 3.84 216.14 ;
		RECT	4.055 216.01 4.105 216.14 ;
		RECT	6.76 216.01 6.81 216.14 ;
		RECT	8.04 216.01 8.09 216.14 ;
		RECT	10.26 216.01 10.31 216.14 ;
		RECT	11.565 216.01 11.615 216.14 ;
		RECT	2.11 216.995 2.16 217.125 ;
		RECT	5.41 216.995 5.46 217.125 ;
		RECT	6.915 216.995 6.965 217.125 ;
		RECT	10.54 216.995 10.59 217.125 ;
		RECT	10.81 216.995 10.86 217.125 ;
		RECT	13.33 216.995 13.38 217.125 ;
		RECT	2.4 217.975 2.45 218.105 ;
		RECT	2.55 217.975 2.6 218.105 ;
		RECT	2.86 217.975 2.91 218.105 ;
		RECT	3.79 217.975 3.84 218.105 ;
		RECT	4.055 217.975 4.105 218.105 ;
		RECT	6.76 217.975 6.81 218.105 ;
		RECT	8.04 217.975 8.09 218.105 ;
		RECT	10.26 217.975 10.31 218.105 ;
		RECT	11.565 217.975 11.615 218.105 ;
		RECT	2.4 218.96 2.45 219.09 ;
		RECT	2.55 218.96 2.6 219.09 ;
		RECT	2.86 218.96 2.91 219.09 ;
		RECT	3.79 218.96 3.84 219.09 ;
		RECT	4.055 218.96 4.105 219.09 ;
		RECT	6.76 218.96 6.81 219.09 ;
		RECT	8.04 218.96 8.09 219.09 ;
		RECT	10.26 218.96 10.31 219.09 ;
		RECT	11.565 218.96 11.615 219.09 ;
		RECT	2.4 219.945 2.45 220.075 ;
		RECT	2.55 219.945 2.6 220.075 ;
		RECT	2.86 219.945 2.91 220.075 ;
		RECT	3.79 219.945 3.84 220.075 ;
		RECT	4.055 219.945 4.105 220.075 ;
		RECT	6.76 219.945 6.81 220.075 ;
		RECT	8.04 219.945 8.09 220.075 ;
		RECT	10.26 219.945 10.31 220.075 ;
		RECT	11.565 219.945 11.615 220.075 ;
		RECT	2.11 220.93 2.16 221.06 ;
		RECT	3.56 220.905 3.69 221.085 ;
		RECT	5.41 220.93 5.46 221.06 ;
		RECT	6.915 220.93 6.965 221.06 ;
		RECT	13.33 220.93 13.38 221.06 ;
		RECT	14.83 220.905 14.96 221.085 ;
		RECT	1.585 222.87 1.715 223.05 ;
		RECT	1.88 222.87 2.01 223.05 ;
		RECT	2.4 222.895 2.45 223.025 ;
		RECT	2.55 222.895 2.6 223.025 ;
		RECT	2.86 222.895 2.91 223.025 ;
		RECT	3.79 222.895 3.84 223.025 ;
		RECT	4.055 222.895 4.105 223.025 ;
		RECT	5.01 222.87 5.14 223.05 ;
		RECT	6.76 222.895 6.81 223.025 ;
		RECT	8.04 222.895 8.09 223.025 ;
		RECT	9.815 222.87 9.945 223.05 ;
		RECT	10.26 222.895 10.31 223.025 ;
		RECT	11.565 222.895 11.615 223.025 ;
		RECT	2.4 223.88 2.45 224.01 ;
		RECT	2.55 223.88 2.6 224.01 ;
		RECT	2.86 223.88 2.91 224.01 ;
		RECT	3.79 223.88 3.84 224.01 ;
		RECT	4.055 223.88 4.105 224.01 ;
		RECT	6.76 223.88 6.81 224.01 ;
		RECT	8.04 223.88 8.09 224.01 ;
		RECT	10.26 223.88 10.31 224.01 ;
		RECT	11.565 223.88 11.615 224.01 ;
		RECT	2.11 224.88 2.16 225.01 ;
		RECT	3.56 224.855 3.69 225.035 ;
		RECT	5.41 224.88 5.46 225.01 ;
		RECT	6.915 224.88 6.965 225.01 ;
		RECT	12.23 224.88 12.28 225.01 ;
		RECT	13.33 224.88 13.38 225.01 ;
		RECT	2.11 225.355 2.16 225.485 ;
		RECT	3.56 225.33 3.69 225.51 ;
		RECT	5.41 225.355 5.46 225.485 ;
		RECT	6.915 225.355 6.965 225.485 ;
		RECT	2.4 225.85 2.45 225.98 ;
		RECT	2.55 225.85 2.6 225.98 ;
		RECT	3.79 225.85 3.84 225.98 ;
		RECT	4.055 225.85 4.105 225.98 ;
		RECT	6.76 225.85 6.81 225.98 ;
		RECT	8.04 225.85 8.09 225.98 ;
		RECT	10.26 225.85 10.31 225.98 ;
		RECT	11.565 225.85 11.615 225.98 ;
		RECT	2.4 226.835 2.45 226.965 ;
		RECT	2.55 226.835 2.6 226.965 ;
		RECT	3.79 226.835 3.84 226.965 ;
		RECT	4.055 226.835 4.105 226.965 ;
		RECT	6.76 226.835 6.81 226.965 ;
		RECT	8.04 226.835 8.09 226.965 ;
		RECT	10.26 226.835 10.31 226.965 ;
		RECT	11.565 226.835 11.615 226.965 ;
		RECT	2.11 227.145 2.16 227.275 ;
		RECT	3.56 227.12 3.69 227.3 ;
		RECT	5.41 227.145 5.46 227.275 ;
		RECT	6.915 227.145 6.965 227.275 ;
		RECT	9.515 227.145 9.565 227.275 ;
		RECT	13.33 227.145 13.38 227.275 ;
		RECT	14.83 227.12 14.96 227.3 ;
		RECT	3.6 228.315 3.65 228.445 ;
		RECT	5.41 228.315 5.46 228.445 ;
		RECT	6.915 228.315 6.965 228.445 ;
		RECT	9.515 228.315 9.565 228.445 ;
		RECT	13.33 228.315 13.38 228.445 ;
		RECT	3.6 187.58 3.65 187.71 ;
		RECT	14.87 187.58 14.92 187.71 ;
		RECT	1.625 187.965 1.675 188.095 ;
		RECT	1.92 187.965 1.97 188.095 ;
		RECT	5.05 187.965 5.1 188.095 ;
		RECT	9.855 187.965 9.905 188.095 ;
		RECT	1.625 188.945 1.675 189.075 ;
		RECT	1.92 188.945 1.97 189.075 ;
		RECT	5.05 188.945 5.1 189.075 ;
		RECT	9.855 188.945 9.905 189.075 ;
		RECT	1.625 190.915 1.675 191.045 ;
		RECT	1.92 190.915 1.97 191.045 ;
		RECT	5.05 190.915 5.1 191.045 ;
		RECT	9.855 190.915 9.905 191.045 ;
		RECT	1.625 191.9 1.675 192.03 ;
		RECT	1.92 191.9 1.97 192.03 ;
		RECT	5.05 191.9 5.1 192.03 ;
		RECT	3.6 193.87 3.65 194 ;
		RECT	14.87 193.87 14.92 194 ;
		RECT	1.625 194.855 1.675 194.985 ;
		RECT	1.92 194.855 1.97 194.985 ;
		RECT	5.05 194.855 5.1 194.985 ;
		RECT	1.625 195.835 1.675 195.965 ;
		RECT	1.92 195.835 1.97 195.965 ;
		RECT	5.05 195.835 5.1 195.965 ;
		RECT	1.625 196.82 1.675 196.95 ;
		RECT	1.92 196.82 1.97 196.95 ;
		RECT	5.05 196.82 5.1 196.95 ;
		RECT	3.6 197.805 3.65 197.935 ;
		RECT	14.87 197.805 14.92 197.935 ;
		RECT	1.625 198.79 1.675 198.92 ;
		RECT	1.92 198.79 1.97 198.92 ;
		RECT	5.05 198.79 5.1 198.92 ;
		RECT	1.585 199.745 1.715 199.925 ;
		RECT	1.88 199.745 2.01 199.925 ;
		RECT	1.625 200.755 1.675 200.885 ;
		RECT	1.92 200.755 1.97 200.885 ;
		RECT	5.05 200.755 5.1 200.885 ;
		RECT	1.625 202.73 1.675 202.86 ;
		RECT	1.92 202.73 1.97 202.86 ;
		RECT	5.05 202.73 5.1 202.86 ;
		RECT	1.625 203.71 1.675 203.84 ;
		RECT	1.92 203.71 1.97 203.84 ;
		RECT	5.05 203.71 5.1 203.84 ;
		RECT	1.625 206.66 1.675 206.79 ;
		RECT	1.92 206.66 1.97 206.79 ;
		RECT	5.05 206.66 5.1 206.79 ;
		RECT	1.625 208.135 1.675 208.265 ;
		RECT	1.92 208.135 1.97 208.265 ;
		RECT	5.05 208.135 5.1 208.265 ;
		RECT	1.625 211.085 1.675 211.215 ;
		RECT	1.92 211.085 1.97 211.215 ;
		RECT	5.05 211.085 5.1 211.215 ;
		RECT	1.625 212.075 1.675 212.205 ;
		RECT	1.92 212.075 1.97 212.205 ;
		RECT	5.05 212.075 5.1 212.205 ;
		RECT	1.625 214.04 1.675 214.17 ;
		RECT	1.92 214.04 1.97 214.17 ;
		RECT	5.05 214.04 5.1 214.17 ;
		RECT	9.83 214.04 9.88 214.17 ;
		RECT	1.585 215 1.715 215.18 ;
		RECT	1.88 215 2.01 215.18 ;
		RECT	1.625 216.01 1.675 216.14 ;
		RECT	1.92 216.01 1.97 216.14 ;
		RECT	5.05 216.01 5.1 216.14 ;
		RECT	9.83 216.01 9.88 216.14 ;
		RECT	3.6 216.995 3.65 217.125 ;
		RECT	14.87 216.995 14.92 217.125 ;
		RECT	1.625 217.975 1.675 218.105 ;
		RECT	1.92 217.975 1.97 218.105 ;
		RECT	5.05 217.975 5.1 218.105 ;
		RECT	9.855 217.975 9.905 218.105 ;
		RECT	1.625 218.96 1.675 219.09 ;
		RECT	1.92 218.96 1.97 219.09 ;
		RECT	5.05 218.96 5.1 219.09 ;
		RECT	9.855 218.96 9.905 219.09 ;
		RECT	1.625 219.945 1.675 220.075 ;
		RECT	1.92 219.945 1.97 220.075 ;
		RECT	5.05 219.945 5.1 220.075 ;
		RECT	9.855 219.945 9.905 220.075 ;
		RECT	1.625 223.88 1.675 224.01 ;
		RECT	1.92 223.88 1.97 224.01 ;
		RECT	5.05 223.88 5.1 224.01 ;
		RECT	9.855 223.88 9.905 224.01 ;
		RECT	1.625 225.85 1.675 225.98 ;
		RECT	1.92 225.85 1.97 225.98 ;
		RECT	5.05 225.85 5.1 225.98 ;
		RECT	9.855 225.85 9.905 225.98 ;
		RECT	0.9 186.645 0.95 186.775 ;
		RECT	1.44 186.645 1.49 186.775 ;
		RECT	3.025 186.645 3.205 186.775 ;
		RECT	4.38 186.645 4.43 186.775 ;
		RECT	6.215 186.645 6.265 186.775 ;
		RECT	6.605 186.645 6.655 186.775 ;
		RECT	7.265 186.645 7.315 186.775 ;
		RECT	8.89 186.645 8.94 186.775 ;
		RECT	9.31 186.645 9.36 186.775 ;
		RECT	12.095 186.645 12.145 186.775 ;
		RECT	12.355 186.645 12.405 186.775 ;
		RECT	13.06 186.645 13.11 186.775 ;
		RECT	14.545 186.645 14.595 186.775 ;
		RECT	0.62 188.455 0.67 188.585 ;
		RECT	1.16 188.455 1.21 188.585 ;
		RECT	4.19 188.455 4.24 188.585 ;
		RECT	7.72 188.455 7.77 188.585 ;
		RECT	14.68 188.455 14.73 188.585 ;
		RECT	0.62 190.46 0.67 190.59 ;
		RECT	1.16 190.46 1.21 190.59 ;
		RECT	4.19 190.46 4.24 190.59 ;
		RECT	7.72 190.46 7.77 190.59 ;
		RECT	14.68 190.46 14.73 190.59 ;
		RECT	0.62 193.375 0.67 193.505 ;
		RECT	1.16 193.375 1.21 193.505 ;
		RECT	4.19 193.375 4.24 193.505 ;
		RECT	7.72 193.375 7.77 193.505 ;
		RECT	14.68 193.375 14.73 193.505 ;
		RECT	0.62 194.36 0.67 194.49 ;
		RECT	1.16 194.36 1.21 194.49 ;
		RECT	4.19 194.36 4.24 194.49 ;
		RECT	7.72 194.36 7.77 194.49 ;
		RECT	14.68 194.36 14.73 194.49 ;
		RECT	0.62 196.33 0.67 196.46 ;
		RECT	1.16 196.33 1.21 196.46 ;
		RECT	4.19 196.33 4.24 196.46 ;
		RECT	7.72 196.33 7.77 196.46 ;
		RECT	14.68 196.33 14.73 196.46 ;
		RECT	0.62 197.31 0.67 197.44 ;
		RECT	1.16 197.31 1.21 197.44 ;
		RECT	4.19 197.31 4.24 197.44 ;
		RECT	7.72 197.31 7.77 197.44 ;
		RECT	14.68 197.31 14.73 197.44 ;
		RECT	0.62 198.295 0.67 198.425 ;
		RECT	1.16 198.295 1.21 198.425 ;
		RECT	4.19 198.295 4.24 198.425 ;
		RECT	7.72 198.295 7.77 198.425 ;
		RECT	14.68 198.295 14.73 198.425 ;
		RECT	0.62 201.25 0.67 201.38 ;
		RECT	1.16 201.25 1.21 201.38 ;
		RECT	4.19 201.25 4.24 201.38 ;
		RECT	7.72 201.25 7.77 201.38 ;
		RECT	14.68 201.25 14.73 201.38 ;
		RECT	0.9 202.235 0.95 202.365 ;
		RECT	1.44 202.235 1.49 202.365 ;
		RECT	3.025 202.235 3.205 202.365 ;
		RECT	6.605 202.235 6.655 202.365 ;
		RECT	7.215 202.235 7.265 202.365 ;
		RECT	12.095 202.235 12.145 202.365 ;
		RECT	12.355 202.235 12.405 202.365 ;
		RECT	13.06 202.235 13.11 202.365 ;
		RECT	14.545 202.235 14.595 202.365 ;
		RECT	0.62 205.185 0.67 205.315 ;
		RECT	1.16 205.185 1.21 205.315 ;
		RECT	4.19 205.185 4.24 205.315 ;
		RECT	7.72 205.185 7.77 205.315 ;
		RECT	14.68 205.185 14.73 205.315 ;
		RECT	0.62 206.17 0.67 206.3 ;
		RECT	1.16 206.17 1.21 206.3 ;
		RECT	4.19 206.17 4.24 206.3 ;
		RECT	7.72 206.17 7.77 206.3 ;
		RECT	14.68 206.17 14.73 206.3 ;
		RECT	8.85 207.44 8.98 207.49 ;
		RECT	9.27 207.44 9.4 207.49 ;
		RECT	10.66 207.44 10.71 207.49 ;
		RECT	12.095 207.44 12.145 207.49 ;
		RECT	12.355 207.44 12.405 207.49 ;
		RECT	13.06 207.44 13.11 207.49 ;
		RECT	0.62 208.63 0.67 208.76 ;
		RECT	1.16 208.63 1.21 208.76 ;
		RECT	4.19 208.63 4.24 208.76 ;
		RECT	7.72 208.63 7.77 208.76 ;
		RECT	13.195 208.63 13.245 208.76 ;
		RECT	14.68 208.63 14.73 208.76 ;
		RECT	0.62 209.61 0.67 209.74 ;
		RECT	1.16 209.61 1.21 209.74 ;
		RECT	4.19 209.61 4.24 209.74 ;
		RECT	7.72 209.61 7.77 209.74 ;
		RECT	14.68 209.61 14.73 209.74 ;
		RECT	0.9 212.565 0.95 212.695 ;
		RECT	1.44 212.565 1.49 212.695 ;
		RECT	3.05 212.54 3.18 212.72 ;
		RECT	4.34 212.54 4.47 212.72 ;
		RECT	6.175 212.54 6.305 212.72 ;
		RECT	6.605 212.565 6.655 212.695 ;
		RECT	7.215 212.565 7.265 212.695 ;
		RECT	8.85 212.54 8.98 212.72 ;
		RECT	9.27 212.54 9.4 212.72 ;
		RECT	12.095 212.565 12.145 212.695 ;
		RECT	12.355 212.565 12.405 212.695 ;
		RECT	13.06 212.565 13.11 212.695 ;
		RECT	14.545 212.565 14.595 212.695 ;
		RECT	0.62 213.55 0.67 213.68 ;
		RECT	1.16 213.55 1.21 213.68 ;
		RECT	4.19 213.55 4.24 213.68 ;
		RECT	7.72 213.55 7.77 213.68 ;
		RECT	14.68 213.55 14.73 213.68 ;
		RECT	0.62 216.5 0.67 216.63 ;
		RECT	1.16 216.5 1.21 216.63 ;
		RECT	4.19 216.5 4.24 216.63 ;
		RECT	7.72 216.5 7.77 216.63 ;
		RECT	14.68 216.5 14.73 216.63 ;
		RECT	0.62 217.485 0.67 217.615 ;
		RECT	1.16 217.485 1.21 217.615 ;
		RECT	4.19 217.485 4.24 217.615 ;
		RECT	7.72 217.485 7.77 217.615 ;
		RECT	14.68 217.485 14.73 217.615 ;
		RECT	0.62 218.47 0.67 218.6 ;
		RECT	1.16 218.47 1.21 218.6 ;
		RECT	4.19 218.47 4.24 218.6 ;
		RECT	7.72 218.47 7.77 218.6 ;
		RECT	14.68 218.47 14.73 218.6 ;
		RECT	0.62 220.435 0.67 220.565 ;
		RECT	1.16 220.435 1.21 220.565 ;
		RECT	4.19 220.435 4.24 220.565 ;
		RECT	7.72 220.435 7.77 220.565 ;
		RECT	14.68 220.435 14.73 220.565 ;
		RECT	0.62 221.215 0.67 221.265 ;
		RECT	1.16 221.215 1.21 221.265 ;
		RECT	0.62 221.42 0.67 221.55 ;
		RECT	1.16 221.42 1.21 221.55 ;
		RECT	4.19 221.42 4.24 221.55 ;
		RECT	7.72 221.42 7.77 221.55 ;
		RECT	14.68 221.42 14.73 221.55 ;
		RECT	0.62 224.34 0.67 224.47 ;
		RECT	1.16 224.34 1.21 224.47 ;
		RECT	4.19 224.34 4.24 224.47 ;
		RECT	7.72 224.34 7.77 224.47 ;
		RECT	14.68 224.34 14.73 224.47 ;
		RECT	0.62 226.34 0.67 226.47 ;
		RECT	1.16 226.34 1.21 226.47 ;
		RECT	4.19 226.34 4.24 226.47 ;
		RECT	7.72 226.34 7.77 226.47 ;
		RECT	14.68 226.34 14.73 226.47 ;
		RECT	0.9 228.085 0.95 228.215 ;
		RECT	1.44 228.085 1.49 228.215 ;
		RECT	3.025 228.085 3.205 228.215 ;
		RECT	4.38 228.085 4.43 228.215 ;
		RECT	6.215 228.085 6.265 228.215 ;
		RECT	6.605 228.085 6.655 228.215 ;
		RECT	7.265 228.085 7.315 228.215 ;
		RECT	8.89 228.085 8.94 228.215 ;
		RECT	9.31 228.085 9.36 228.215 ;
		RECT	12.095 228.085 12.145 228.215 ;
		RECT	12.355 228.085 12.405 228.215 ;
		RECT	13.06 228.085 13.11 228.215 ;
		RECT	14.545 228.085 14.595 228.215 ;
		RECT	4.38 202.235 4.43 202.365 ;
		RECT	6.215 202.235 6.265 202.365 ;
		RECT	8.89 202.235 8.94 202.365 ;
		RECT	9.31 202.235 9.36 202.365 ;
		RECT	2.11 186.875 2.16 187.005 ;
		RECT	3.6 186.875 3.65 187.005 ;
		RECT	5.41 186.875 5.46 187.005 ;
		RECT	13.33 186.875 13.38 187.005 ;
		RECT	14.87 186.875 14.92 187.005 ;
		RECT	2.72 187.965 2.77 188.095 ;
		RECT	9.1 187.965 9.15 188.095 ;
		RECT	10.81 187.965 10.86 188.095 ;
		RECT	2.72 188.945 2.77 189.075 ;
		RECT	9.1 188.945 9.15 189.075 ;
		RECT	10.81 188.945 10.86 189.075 ;
		RECT	2.72 190.915 2.77 191.045 ;
		RECT	9.1 190.915 9.15 191.045 ;
		RECT	10.81 190.915 10.86 191.045 ;
		RECT	2.72 191.9 2.77 192.03 ;
		RECT	9.1 191.9 9.15 192.03 ;
		RECT	10.81 191.9 10.86 192.03 ;
		RECT	2.11 192.885 2.16 193.015 ;
		RECT	5.41 192.885 5.46 193.015 ;
		RECT	6.44 192.885 6.49 193.015 ;
		RECT	13.33 192.885 13.38 193.015 ;
		RECT	2.72 194.855 2.77 194.985 ;
		RECT	9.1 194.855 9.15 194.985 ;
		RECT	2.72 195.835 2.77 195.965 ;
		RECT	9.1 195.835 9.15 195.965 ;
		RECT	2.72 196.82 2.77 196.95 ;
		RECT	9.1 196.82 9.15 196.95 ;
		RECT	2.72 198.79 2.77 198.92 ;
		RECT	9.1 198.79 9.15 198.92 ;
		RECT	2.72 199.77 2.77 199.9 ;
		RECT	9.1 199.77 9.15 199.9 ;
		RECT	2.72 200.755 2.77 200.885 ;
		RECT	9.1 200.755 9.15 200.885 ;
		RECT	2.72 202.73 2.77 202.86 ;
		RECT	9.1 202.73 9.15 202.86 ;
		RECT	2.72 203.71 2.77 203.84 ;
		RECT	9.1 203.71 9.15 203.84 ;
		RECT	2.72 206.66 2.77 206.79 ;
		RECT	9.1 206.66 9.15 206.79 ;
		RECT	2.72 208.135 2.77 208.265 ;
		RECT	9.1 208.135 9.15 208.265 ;
		RECT	2.72 211.085 2.77 211.215 ;
		RECT	9.1 211.085 9.15 211.215 ;
		RECT	2.72 212.075 2.77 212.205 ;
		RECT	9.1 212.075 9.15 212.205 ;
		RECT	2.72 214.04 2.77 214.17 ;
		RECT	9.1 214.04 9.15 214.17 ;
		RECT	2.72 215.025 2.77 215.155 ;
		RECT	9.1 215.025 9.15 215.155 ;
		RECT	2.72 216.01 2.77 216.14 ;
		RECT	9.1 216.01 9.15 216.14 ;
		RECT	2.72 217.975 2.77 218.105 ;
		RECT	9.1 217.975 9.15 218.105 ;
		RECT	2.72 218.96 2.77 219.09 ;
		RECT	9.1 218.96 9.15 219.09 ;
		RECT	2.72 219.945 2.77 220.075 ;
		RECT	9.1 219.945 9.15 220.075 ;
		RECT	2.11 221.915 2.16 222.045 ;
		RECT	3.56 221.89 3.69 222.07 ;
		RECT	5.41 221.915 5.46 222.045 ;
		RECT	6.915 221.915 6.965 222.045 ;
		RECT	13.33 221.915 13.38 222.045 ;
		RECT	14.83 221.89 14.96 222.07 ;
		RECT	2.72 222.895 2.77 223.025 ;
		RECT	9.1 222.895 9.15 223.025 ;
		RECT	10.81 222.895 10.86 223.025 ;
		RECT	2.72 223.88 2.77 224.01 ;
		RECT	9.1 223.88 9.15 224.01 ;
		RECT	10.81 223.88 10.86 224.01 ;
		RECT	2.72 225.85 2.77 225.98 ;
		RECT	9.1 225.85 9.15 225.98 ;
		RECT	10.81 225.85 10.86 225.98 ;
		RECT	2.72 226.835 2.77 226.965 ;
		RECT	9.1 226.835 9.15 226.965 ;
		RECT	10.81 226.835 10.86 226.965 ;
		RECT	3.6 227.855 3.65 227.985 ;
		RECT	5.41 227.855 5.46 227.985 ;
		RECT	6.915 227.855 6.965 227.985 ;
		RECT	9.515 227.855 9.565 227.985 ;
		RECT	13.33 227.855 13.38 227.985 ;
		RECT	14.87 227.855 14.92 227.985 ;
		RECT	3.6 192.885 3.65 193.015 ;
		RECT	14.87 192.885 14.92 193.015 ;
		RECT	21.685 0.425 21.865 0.555 ;
		RECT	15.775 0.655 15.825 0.785 ;
		RECT	20.295 0.655 20.345 0.785 ;
		RECT	15.575 0.655 15.625 0.785 ;
		RECT	20.495 0.655 20.545 0.785 ;
		RECT	21.51 0.425 21.56 0.555 ;
		RECT	21.685 414.305 21.865 414.435 ;
		RECT	15.775 414.075 15.825 414.205 ;
		RECT	20.295 414.075 20.345 414.205 ;
		RECT	15.575 414.075 15.625 414.205 ;
		RECT	20.495 414.075 20.545 414.205 ;
		RECT	21.51 414.305 21.56 414.435 ;
		RECT	15.375 3.305 15.425 3.435 ;
		RECT	20.695 3.305 20.745 3.435 ;
		RECT	15.575 3.535 15.625 3.665 ;
		RECT	15.575 1.115 15.625 1.245 ;
		RECT	20.495 3.535 20.545 3.665 ;
		RECT	20.495 1.115 20.545 1.245 ;
		RECT	15.775 3.535 15.825 3.665 ;
		RECT	15.775 1.115 15.825 1.245 ;
		RECT	20.295 3.535 20.345 3.665 ;
		RECT	20.295 1.115 20.345 1.245 ;
		RECT	15.375 184.745 15.425 184.875 ;
		RECT	20.695 184.745 20.745 184.875 ;
		RECT	15.575 184.975 15.625 185.105 ;
		RECT	15.575 182.555 15.625 182.685 ;
		RECT	20.495 184.975 20.545 185.105 ;
		RECT	20.495 182.555 20.545 182.685 ;
		RECT	15.775 184.975 15.825 185.105 ;
		RECT	15.775 182.555 15.825 182.685 ;
		RECT	20.295 184.975 20.345 185.105 ;
		RECT	20.295 182.555 20.345 182.685 ;
		RECT	15.375 181.865 15.425 181.995 ;
		RECT	20.695 181.865 20.745 181.995 ;
		RECT	15.575 182.095 15.625 182.225 ;
		RECT	15.575 179.675 15.625 179.805 ;
		RECT	20.495 182.095 20.545 182.225 ;
		RECT	20.495 179.675 20.545 179.805 ;
		RECT	15.775 182.095 15.825 182.225 ;
		RECT	15.775 179.675 15.825 179.805 ;
		RECT	20.295 182.095 20.345 182.225 ;
		RECT	20.295 179.675 20.345 179.805 ;
		RECT	15.375 155.945 15.425 156.075 ;
		RECT	20.695 155.945 20.745 156.075 ;
		RECT	15.575 156.175 15.625 156.305 ;
		RECT	15.575 153.755 15.625 153.885 ;
		RECT	20.495 156.175 20.545 156.305 ;
		RECT	20.495 153.755 20.545 153.885 ;
		RECT	15.775 156.175 15.825 156.305 ;
		RECT	15.775 153.755 15.825 153.885 ;
		RECT	20.295 156.175 20.345 156.305 ;
		RECT	20.295 153.755 20.345 153.885 ;
		RECT	15.375 153.065 15.425 153.195 ;
		RECT	20.695 153.065 20.745 153.195 ;
		RECT	15.575 153.295 15.625 153.425 ;
		RECT	15.575 150.875 15.625 151.005 ;
		RECT	20.495 153.295 20.545 153.425 ;
		RECT	20.495 150.875 20.545 151.005 ;
		RECT	15.775 153.295 15.825 153.425 ;
		RECT	15.775 150.875 15.825 151.005 ;
		RECT	20.295 153.295 20.345 153.425 ;
		RECT	20.295 150.875 20.345 151.005 ;
		RECT	15.375 150.185 15.425 150.315 ;
		RECT	20.695 150.185 20.745 150.315 ;
		RECT	15.575 150.415 15.625 150.545 ;
		RECT	15.575 147.995 15.625 148.125 ;
		RECT	20.495 150.415 20.545 150.545 ;
		RECT	20.495 147.995 20.545 148.125 ;
		RECT	15.775 150.415 15.825 150.545 ;
		RECT	15.775 147.995 15.825 148.125 ;
		RECT	20.295 150.415 20.345 150.545 ;
		RECT	20.295 147.995 20.345 148.125 ;
		RECT	15.375 147.305 15.425 147.435 ;
		RECT	20.695 147.305 20.745 147.435 ;
		RECT	15.575 147.535 15.625 147.665 ;
		RECT	15.575 145.115 15.625 145.245 ;
		RECT	20.495 147.535 20.545 147.665 ;
		RECT	20.495 145.115 20.545 145.245 ;
		RECT	15.775 147.535 15.825 147.665 ;
		RECT	15.775 145.115 15.825 145.245 ;
		RECT	20.295 147.535 20.345 147.665 ;
		RECT	20.295 145.115 20.345 145.245 ;
		RECT	15.375 144.425 15.425 144.555 ;
		RECT	20.695 144.425 20.745 144.555 ;
		RECT	15.575 144.655 15.625 144.785 ;
		RECT	15.575 142.235 15.625 142.365 ;
		RECT	20.495 144.655 20.545 144.785 ;
		RECT	20.495 142.235 20.545 142.365 ;
		RECT	15.775 144.655 15.825 144.785 ;
		RECT	15.775 142.235 15.825 142.365 ;
		RECT	20.295 144.655 20.345 144.785 ;
		RECT	20.295 142.235 20.345 142.365 ;
		RECT	15.375 141.545 15.425 141.675 ;
		RECT	20.695 141.545 20.745 141.675 ;
		RECT	15.575 141.775 15.625 141.905 ;
		RECT	15.575 139.355 15.625 139.485 ;
		RECT	20.495 141.775 20.545 141.905 ;
		RECT	20.495 139.355 20.545 139.485 ;
		RECT	15.775 141.775 15.825 141.905 ;
		RECT	15.775 139.355 15.825 139.485 ;
		RECT	20.295 141.775 20.345 141.905 ;
		RECT	20.295 139.355 20.345 139.485 ;
		RECT	15.375 138.665 15.425 138.795 ;
		RECT	20.695 138.665 20.745 138.795 ;
		RECT	15.575 138.895 15.625 139.025 ;
		RECT	15.575 136.475 15.625 136.605 ;
		RECT	20.495 138.895 20.545 139.025 ;
		RECT	20.495 136.475 20.545 136.605 ;
		RECT	15.775 138.895 15.825 139.025 ;
		RECT	15.775 136.475 15.825 136.605 ;
		RECT	20.295 138.895 20.345 139.025 ;
		RECT	20.295 136.475 20.345 136.605 ;
		RECT	15.375 135.785 15.425 135.915 ;
		RECT	20.695 135.785 20.745 135.915 ;
		RECT	15.575 136.015 15.625 136.145 ;
		RECT	15.575 133.595 15.625 133.725 ;
		RECT	20.495 136.015 20.545 136.145 ;
		RECT	20.495 133.595 20.545 133.725 ;
		RECT	15.775 136.015 15.825 136.145 ;
		RECT	15.775 133.595 15.825 133.725 ;
		RECT	20.295 136.015 20.345 136.145 ;
		RECT	20.295 133.595 20.345 133.725 ;
		RECT	15.375 132.905 15.425 133.035 ;
		RECT	20.695 132.905 20.745 133.035 ;
		RECT	15.575 133.135 15.625 133.265 ;
		RECT	15.575 130.715 15.625 130.845 ;
		RECT	20.495 133.135 20.545 133.265 ;
		RECT	20.495 130.715 20.545 130.845 ;
		RECT	15.775 133.135 15.825 133.265 ;
		RECT	15.775 130.715 15.825 130.845 ;
		RECT	20.295 133.135 20.345 133.265 ;
		RECT	20.295 130.715 20.345 130.845 ;
		RECT	15.375 130.025 15.425 130.155 ;
		RECT	20.695 130.025 20.745 130.155 ;
		RECT	15.575 130.255 15.625 130.385 ;
		RECT	15.575 127.835 15.625 127.965 ;
		RECT	20.495 130.255 20.545 130.385 ;
		RECT	20.495 127.835 20.545 127.965 ;
		RECT	15.775 130.255 15.825 130.385 ;
		RECT	15.775 127.835 15.825 127.965 ;
		RECT	20.295 130.255 20.345 130.385 ;
		RECT	20.295 127.835 20.345 127.965 ;
		RECT	15.375 178.985 15.425 179.115 ;
		RECT	20.695 178.985 20.745 179.115 ;
		RECT	15.575 179.215 15.625 179.345 ;
		RECT	15.575 176.795 15.625 176.925 ;
		RECT	20.495 179.215 20.545 179.345 ;
		RECT	20.495 176.795 20.545 176.925 ;
		RECT	15.775 179.215 15.825 179.345 ;
		RECT	15.775 176.795 15.825 176.925 ;
		RECT	20.295 179.215 20.345 179.345 ;
		RECT	20.295 176.795 20.345 176.925 ;
		RECT	15.375 127.145 15.425 127.275 ;
		RECT	20.695 127.145 20.745 127.275 ;
		RECT	15.575 127.375 15.625 127.505 ;
		RECT	15.575 124.955 15.625 125.085 ;
		RECT	20.495 127.375 20.545 127.505 ;
		RECT	20.495 124.955 20.545 125.085 ;
		RECT	15.775 127.375 15.825 127.505 ;
		RECT	15.775 124.955 15.825 125.085 ;
		RECT	20.295 127.375 20.345 127.505 ;
		RECT	20.295 124.955 20.345 125.085 ;
		RECT	15.375 124.265 15.425 124.395 ;
		RECT	20.695 124.265 20.745 124.395 ;
		RECT	15.575 124.495 15.625 124.625 ;
		RECT	15.575 122.075 15.625 122.205 ;
		RECT	20.495 124.495 20.545 124.625 ;
		RECT	20.495 122.075 20.545 122.205 ;
		RECT	15.775 124.495 15.825 124.625 ;
		RECT	15.775 122.075 15.825 122.205 ;
		RECT	20.295 124.495 20.345 124.625 ;
		RECT	20.295 122.075 20.345 122.205 ;
		RECT	15.375 121.385 15.425 121.515 ;
		RECT	20.695 121.385 20.745 121.515 ;
		RECT	15.575 121.615 15.625 121.745 ;
		RECT	15.575 119.195 15.625 119.325 ;
		RECT	20.495 121.615 20.545 121.745 ;
		RECT	20.495 119.195 20.545 119.325 ;
		RECT	15.775 121.615 15.825 121.745 ;
		RECT	15.775 119.195 15.825 119.325 ;
		RECT	20.295 121.615 20.345 121.745 ;
		RECT	20.295 119.195 20.345 119.325 ;
		RECT	15.375 118.505 15.425 118.635 ;
		RECT	20.695 118.505 20.745 118.635 ;
		RECT	15.575 118.735 15.625 118.865 ;
		RECT	15.575 116.315 15.625 116.445 ;
		RECT	20.495 118.735 20.545 118.865 ;
		RECT	20.495 116.315 20.545 116.445 ;
		RECT	15.775 118.735 15.825 118.865 ;
		RECT	15.775 116.315 15.825 116.445 ;
		RECT	20.295 118.735 20.345 118.865 ;
		RECT	20.295 116.315 20.345 116.445 ;
		RECT	15.375 115.625 15.425 115.755 ;
		RECT	20.695 115.625 20.745 115.755 ;
		RECT	15.575 115.855 15.625 115.985 ;
		RECT	15.575 113.435 15.625 113.565 ;
		RECT	20.495 115.855 20.545 115.985 ;
		RECT	20.495 113.435 20.545 113.565 ;
		RECT	15.775 115.855 15.825 115.985 ;
		RECT	15.775 113.435 15.825 113.565 ;
		RECT	20.295 115.855 20.345 115.985 ;
		RECT	20.295 113.435 20.345 113.565 ;
		RECT	15.375 112.745 15.425 112.875 ;
		RECT	20.695 112.745 20.745 112.875 ;
		RECT	15.575 112.975 15.625 113.105 ;
		RECT	15.575 110.555 15.625 110.685 ;
		RECT	20.495 112.975 20.545 113.105 ;
		RECT	20.495 110.555 20.545 110.685 ;
		RECT	15.775 112.975 15.825 113.105 ;
		RECT	15.775 110.555 15.825 110.685 ;
		RECT	20.295 112.975 20.345 113.105 ;
		RECT	20.295 110.555 20.345 110.685 ;
		RECT	15.375 109.865 15.425 109.995 ;
		RECT	20.695 109.865 20.745 109.995 ;
		RECT	15.575 110.095 15.625 110.225 ;
		RECT	15.575 107.675 15.625 107.805 ;
		RECT	20.495 110.095 20.545 110.225 ;
		RECT	20.495 107.675 20.545 107.805 ;
		RECT	15.775 110.095 15.825 110.225 ;
		RECT	15.775 107.675 15.825 107.805 ;
		RECT	20.295 110.095 20.345 110.225 ;
		RECT	20.295 107.675 20.345 107.805 ;
		RECT	15.375 106.985 15.425 107.115 ;
		RECT	20.695 106.985 20.745 107.115 ;
		RECT	15.575 107.215 15.625 107.345 ;
		RECT	15.575 104.795 15.625 104.925 ;
		RECT	20.495 107.215 20.545 107.345 ;
		RECT	20.495 104.795 20.545 104.925 ;
		RECT	15.775 107.215 15.825 107.345 ;
		RECT	15.775 104.795 15.825 104.925 ;
		RECT	20.295 107.215 20.345 107.345 ;
		RECT	20.295 104.795 20.345 104.925 ;
		RECT	15.375 104.105 15.425 104.235 ;
		RECT	20.695 104.105 20.745 104.235 ;
		RECT	15.575 104.335 15.625 104.465 ;
		RECT	15.575 101.915 15.625 102.045 ;
		RECT	20.495 104.335 20.545 104.465 ;
		RECT	20.495 101.915 20.545 102.045 ;
		RECT	15.775 104.335 15.825 104.465 ;
		RECT	15.775 101.915 15.825 102.045 ;
		RECT	20.295 104.335 20.345 104.465 ;
		RECT	20.295 101.915 20.345 102.045 ;
		RECT	15.375 101.225 15.425 101.355 ;
		RECT	20.695 101.225 20.745 101.355 ;
		RECT	15.575 101.455 15.625 101.585 ;
		RECT	15.575 99.035 15.625 99.165 ;
		RECT	20.495 101.455 20.545 101.585 ;
		RECT	20.495 99.035 20.545 99.165 ;
		RECT	15.775 101.455 15.825 101.585 ;
		RECT	15.775 99.035 15.825 99.165 ;
		RECT	20.295 101.455 20.345 101.585 ;
		RECT	20.295 99.035 20.345 99.165 ;
		RECT	15.375 176.105 15.425 176.235 ;
		RECT	20.695 176.105 20.745 176.235 ;
		RECT	15.575 176.335 15.625 176.465 ;
		RECT	15.575 173.915 15.625 174.045 ;
		RECT	20.495 176.335 20.545 176.465 ;
		RECT	20.495 173.915 20.545 174.045 ;
		RECT	15.775 176.335 15.825 176.465 ;
		RECT	15.775 173.915 15.825 174.045 ;
		RECT	20.295 176.335 20.345 176.465 ;
		RECT	20.295 173.915 20.345 174.045 ;
		RECT	15.375 98.345 15.425 98.475 ;
		RECT	20.695 98.345 20.745 98.475 ;
		RECT	15.575 98.575 15.625 98.705 ;
		RECT	15.575 96.155 15.625 96.285 ;
		RECT	20.495 98.575 20.545 98.705 ;
		RECT	20.495 96.155 20.545 96.285 ;
		RECT	15.775 98.575 15.825 98.705 ;
		RECT	15.775 96.155 15.825 96.285 ;
		RECT	20.295 98.575 20.345 98.705 ;
		RECT	20.295 96.155 20.345 96.285 ;
		RECT	15.375 95.465 15.425 95.595 ;
		RECT	20.695 95.465 20.745 95.595 ;
		RECT	15.575 95.695 15.625 95.825 ;
		RECT	15.575 93.275 15.625 93.405 ;
		RECT	20.495 95.695 20.545 95.825 ;
		RECT	20.495 93.275 20.545 93.405 ;
		RECT	15.775 95.695 15.825 95.825 ;
		RECT	15.775 93.275 15.825 93.405 ;
		RECT	20.295 95.695 20.345 95.825 ;
		RECT	20.295 93.275 20.345 93.405 ;
		RECT	15.375 92.585 15.425 92.715 ;
		RECT	20.695 92.585 20.745 92.715 ;
		RECT	15.575 92.815 15.625 92.945 ;
		RECT	15.575 90.395 15.625 90.525 ;
		RECT	20.495 92.815 20.545 92.945 ;
		RECT	20.495 90.395 20.545 90.525 ;
		RECT	15.775 92.815 15.825 92.945 ;
		RECT	15.775 90.395 15.825 90.525 ;
		RECT	20.295 92.815 20.345 92.945 ;
		RECT	20.295 90.395 20.345 90.525 ;
		RECT	15.375 89.705 15.425 89.835 ;
		RECT	20.695 89.705 20.745 89.835 ;
		RECT	15.575 89.935 15.625 90.065 ;
		RECT	15.575 87.515 15.625 87.645 ;
		RECT	20.495 89.935 20.545 90.065 ;
		RECT	20.495 87.515 20.545 87.645 ;
		RECT	15.775 89.935 15.825 90.065 ;
		RECT	15.775 87.515 15.825 87.645 ;
		RECT	20.295 89.935 20.345 90.065 ;
		RECT	20.295 87.515 20.345 87.645 ;
		RECT	15.375 86.825 15.425 86.955 ;
		RECT	20.695 86.825 20.745 86.955 ;
		RECT	15.575 87.055 15.625 87.185 ;
		RECT	15.575 84.635 15.625 84.765 ;
		RECT	20.495 87.055 20.545 87.185 ;
		RECT	20.495 84.635 20.545 84.765 ;
		RECT	15.775 87.055 15.825 87.185 ;
		RECT	15.775 84.635 15.825 84.765 ;
		RECT	20.295 87.055 20.345 87.185 ;
		RECT	20.295 84.635 20.345 84.765 ;
		RECT	15.375 83.945 15.425 84.075 ;
		RECT	20.695 83.945 20.745 84.075 ;
		RECT	15.575 84.175 15.625 84.305 ;
		RECT	15.575 81.755 15.625 81.885 ;
		RECT	20.495 84.175 20.545 84.305 ;
		RECT	20.495 81.755 20.545 81.885 ;
		RECT	15.775 84.175 15.825 84.305 ;
		RECT	15.775 81.755 15.825 81.885 ;
		RECT	20.295 84.175 20.345 84.305 ;
		RECT	20.295 81.755 20.345 81.885 ;
		RECT	15.375 81.065 15.425 81.195 ;
		RECT	20.695 81.065 20.745 81.195 ;
		RECT	15.575 81.295 15.625 81.425 ;
		RECT	15.575 78.875 15.625 79.005 ;
		RECT	20.495 81.295 20.545 81.425 ;
		RECT	20.495 78.875 20.545 79.005 ;
		RECT	15.775 81.295 15.825 81.425 ;
		RECT	15.775 78.875 15.825 79.005 ;
		RECT	20.295 81.295 20.345 81.425 ;
		RECT	20.295 78.875 20.345 79.005 ;
		RECT	15.375 78.185 15.425 78.315 ;
		RECT	20.695 78.185 20.745 78.315 ;
		RECT	15.575 78.415 15.625 78.545 ;
		RECT	15.575 75.995 15.625 76.125 ;
		RECT	20.495 78.415 20.545 78.545 ;
		RECT	20.495 75.995 20.545 76.125 ;
		RECT	15.775 78.415 15.825 78.545 ;
		RECT	15.775 75.995 15.825 76.125 ;
		RECT	20.295 78.415 20.345 78.545 ;
		RECT	20.295 75.995 20.345 76.125 ;
		RECT	15.375 75.305 15.425 75.435 ;
		RECT	20.695 75.305 20.745 75.435 ;
		RECT	15.575 75.535 15.625 75.665 ;
		RECT	15.575 73.115 15.625 73.245 ;
		RECT	20.495 75.535 20.545 75.665 ;
		RECT	20.495 73.115 20.545 73.245 ;
		RECT	15.775 75.535 15.825 75.665 ;
		RECT	15.775 73.115 15.825 73.245 ;
		RECT	20.295 75.535 20.345 75.665 ;
		RECT	20.295 73.115 20.345 73.245 ;
		RECT	15.375 72.425 15.425 72.555 ;
		RECT	20.695 72.425 20.745 72.555 ;
		RECT	15.575 72.655 15.625 72.785 ;
		RECT	15.575 70.235 15.625 70.365 ;
		RECT	20.495 72.655 20.545 72.785 ;
		RECT	20.495 70.235 20.545 70.365 ;
		RECT	15.775 72.655 15.825 72.785 ;
		RECT	15.775 70.235 15.825 70.365 ;
		RECT	20.295 72.655 20.345 72.785 ;
		RECT	20.295 70.235 20.345 70.365 ;
		RECT	15.375 173.225 15.425 173.355 ;
		RECT	20.695 173.225 20.745 173.355 ;
		RECT	15.575 173.455 15.625 173.585 ;
		RECT	15.575 171.035 15.625 171.165 ;
		RECT	20.495 173.455 20.545 173.585 ;
		RECT	20.495 171.035 20.545 171.165 ;
		RECT	15.775 173.455 15.825 173.585 ;
		RECT	15.775 171.035 15.825 171.165 ;
		RECT	20.295 173.455 20.345 173.585 ;
		RECT	20.295 171.035 20.345 171.165 ;
		RECT	15.375 69.545 15.425 69.675 ;
		RECT	20.695 69.545 20.745 69.675 ;
		RECT	15.575 69.775 15.625 69.905 ;
		RECT	15.575 67.355 15.625 67.485 ;
		RECT	20.495 69.775 20.545 69.905 ;
		RECT	20.495 67.355 20.545 67.485 ;
		RECT	15.775 69.775 15.825 69.905 ;
		RECT	15.775 67.355 15.825 67.485 ;
		RECT	20.295 69.775 20.345 69.905 ;
		RECT	20.295 67.355 20.345 67.485 ;
		RECT	15.375 66.665 15.425 66.795 ;
		RECT	20.695 66.665 20.745 66.795 ;
		RECT	15.575 66.895 15.625 67.025 ;
		RECT	15.575 64.475 15.625 64.605 ;
		RECT	20.495 66.895 20.545 67.025 ;
		RECT	20.495 64.475 20.545 64.605 ;
		RECT	15.775 66.895 15.825 67.025 ;
		RECT	15.775 64.475 15.825 64.605 ;
		RECT	20.295 66.895 20.345 67.025 ;
		RECT	20.295 64.475 20.345 64.605 ;
		RECT	15.375 63.785 15.425 63.915 ;
		RECT	20.695 63.785 20.745 63.915 ;
		RECT	15.575 64.015 15.625 64.145 ;
		RECT	15.575 61.595 15.625 61.725 ;
		RECT	20.495 64.015 20.545 64.145 ;
		RECT	20.495 61.595 20.545 61.725 ;
		RECT	15.775 64.015 15.825 64.145 ;
		RECT	15.775 61.595 15.825 61.725 ;
		RECT	20.295 64.015 20.345 64.145 ;
		RECT	20.295 61.595 20.345 61.725 ;
		RECT	15.375 60.905 15.425 61.035 ;
		RECT	20.695 60.905 20.745 61.035 ;
		RECT	15.575 61.135 15.625 61.265 ;
		RECT	15.575 58.715 15.625 58.845 ;
		RECT	20.495 61.135 20.545 61.265 ;
		RECT	20.495 58.715 20.545 58.845 ;
		RECT	15.775 61.135 15.825 61.265 ;
		RECT	15.775 58.715 15.825 58.845 ;
		RECT	20.295 61.135 20.345 61.265 ;
		RECT	20.295 58.715 20.345 58.845 ;
		RECT	15.375 58.025 15.425 58.155 ;
		RECT	20.695 58.025 20.745 58.155 ;
		RECT	15.575 58.255 15.625 58.385 ;
		RECT	15.575 55.835 15.625 55.965 ;
		RECT	20.495 58.255 20.545 58.385 ;
		RECT	20.495 55.835 20.545 55.965 ;
		RECT	15.775 58.255 15.825 58.385 ;
		RECT	15.775 55.835 15.825 55.965 ;
		RECT	20.295 58.255 20.345 58.385 ;
		RECT	20.295 55.835 20.345 55.965 ;
		RECT	15.375 55.145 15.425 55.275 ;
		RECT	20.695 55.145 20.745 55.275 ;
		RECT	15.575 55.375 15.625 55.505 ;
		RECT	15.575 52.955 15.625 53.085 ;
		RECT	20.495 55.375 20.545 55.505 ;
		RECT	20.495 52.955 20.545 53.085 ;
		RECT	15.775 55.375 15.825 55.505 ;
		RECT	15.775 52.955 15.825 53.085 ;
		RECT	20.295 55.375 20.345 55.505 ;
		RECT	20.295 52.955 20.345 53.085 ;
		RECT	15.375 52.265 15.425 52.395 ;
		RECT	20.695 52.265 20.745 52.395 ;
		RECT	15.575 52.495 15.625 52.625 ;
		RECT	15.575 50.075 15.625 50.205 ;
		RECT	20.495 52.495 20.545 52.625 ;
		RECT	20.495 50.075 20.545 50.205 ;
		RECT	15.775 52.495 15.825 52.625 ;
		RECT	15.775 50.075 15.825 50.205 ;
		RECT	20.295 52.495 20.345 52.625 ;
		RECT	20.295 50.075 20.345 50.205 ;
		RECT	15.375 49.385 15.425 49.515 ;
		RECT	20.695 49.385 20.745 49.515 ;
		RECT	15.575 49.615 15.625 49.745 ;
		RECT	15.575 47.195 15.625 47.325 ;
		RECT	20.495 49.615 20.545 49.745 ;
		RECT	20.495 47.195 20.545 47.325 ;
		RECT	15.775 49.615 15.825 49.745 ;
		RECT	15.775 47.195 15.825 47.325 ;
		RECT	20.295 49.615 20.345 49.745 ;
		RECT	20.295 47.195 20.345 47.325 ;
		RECT	15.375 46.505 15.425 46.635 ;
		RECT	20.695 46.505 20.745 46.635 ;
		RECT	15.575 46.735 15.625 46.865 ;
		RECT	15.575 44.315 15.625 44.445 ;
		RECT	20.495 46.735 20.545 46.865 ;
		RECT	20.495 44.315 20.545 44.445 ;
		RECT	15.775 46.735 15.825 46.865 ;
		RECT	15.775 44.315 15.825 44.445 ;
		RECT	20.295 46.735 20.345 46.865 ;
		RECT	20.295 44.315 20.345 44.445 ;
		RECT	15.375 43.625 15.425 43.755 ;
		RECT	20.695 43.625 20.745 43.755 ;
		RECT	15.575 43.855 15.625 43.985 ;
		RECT	15.575 41.435 15.625 41.565 ;
		RECT	20.495 43.855 20.545 43.985 ;
		RECT	20.495 41.435 20.545 41.565 ;
		RECT	15.775 43.855 15.825 43.985 ;
		RECT	15.775 41.435 15.825 41.565 ;
		RECT	20.295 43.855 20.345 43.985 ;
		RECT	20.295 41.435 20.345 41.565 ;
		RECT	15.375 170.345 15.425 170.475 ;
		RECT	20.695 170.345 20.745 170.475 ;
		RECT	15.575 170.575 15.625 170.705 ;
		RECT	15.575 168.155 15.625 168.285 ;
		RECT	20.495 170.575 20.545 170.705 ;
		RECT	20.495 168.155 20.545 168.285 ;
		RECT	15.775 170.575 15.825 170.705 ;
		RECT	15.775 168.155 15.825 168.285 ;
		RECT	20.295 170.575 20.345 170.705 ;
		RECT	20.295 168.155 20.345 168.285 ;
		RECT	15.375 40.745 15.425 40.875 ;
		RECT	20.695 40.745 20.745 40.875 ;
		RECT	15.575 40.975 15.625 41.105 ;
		RECT	15.575 38.555 15.625 38.685 ;
		RECT	20.495 40.975 20.545 41.105 ;
		RECT	20.495 38.555 20.545 38.685 ;
		RECT	15.775 40.975 15.825 41.105 ;
		RECT	15.775 38.555 15.825 38.685 ;
		RECT	20.295 40.975 20.345 41.105 ;
		RECT	20.295 38.555 20.345 38.685 ;
		RECT	15.375 37.865 15.425 37.995 ;
		RECT	20.695 37.865 20.745 37.995 ;
		RECT	15.575 38.095 15.625 38.225 ;
		RECT	15.575 35.675 15.625 35.805 ;
		RECT	20.495 38.095 20.545 38.225 ;
		RECT	20.495 35.675 20.545 35.805 ;
		RECT	15.775 38.095 15.825 38.225 ;
		RECT	15.775 35.675 15.825 35.805 ;
		RECT	20.295 38.095 20.345 38.225 ;
		RECT	20.295 35.675 20.345 35.805 ;
		RECT	15.375 34.985 15.425 35.115 ;
		RECT	20.695 34.985 20.745 35.115 ;
		RECT	15.575 35.215 15.625 35.345 ;
		RECT	15.575 32.795 15.625 32.925 ;
		RECT	20.495 35.215 20.545 35.345 ;
		RECT	20.495 32.795 20.545 32.925 ;
		RECT	15.775 35.215 15.825 35.345 ;
		RECT	15.775 32.795 15.825 32.925 ;
		RECT	20.295 35.215 20.345 35.345 ;
		RECT	20.295 32.795 20.345 32.925 ;
		RECT	15.375 32.105 15.425 32.235 ;
		RECT	20.695 32.105 20.745 32.235 ;
		RECT	15.575 32.335 15.625 32.465 ;
		RECT	15.575 29.915 15.625 30.045 ;
		RECT	20.495 32.335 20.545 32.465 ;
		RECT	20.495 29.915 20.545 30.045 ;
		RECT	15.775 32.335 15.825 32.465 ;
		RECT	15.775 29.915 15.825 30.045 ;
		RECT	20.295 32.335 20.345 32.465 ;
		RECT	20.295 29.915 20.345 30.045 ;
		RECT	15.375 29.225 15.425 29.355 ;
		RECT	20.695 29.225 20.745 29.355 ;
		RECT	15.575 29.455 15.625 29.585 ;
		RECT	15.575 27.035 15.625 27.165 ;
		RECT	20.495 29.455 20.545 29.585 ;
		RECT	20.495 27.035 20.545 27.165 ;
		RECT	15.775 29.455 15.825 29.585 ;
		RECT	15.775 27.035 15.825 27.165 ;
		RECT	20.295 29.455 20.345 29.585 ;
		RECT	20.295 27.035 20.345 27.165 ;
		RECT	15.375 26.345 15.425 26.475 ;
		RECT	20.695 26.345 20.745 26.475 ;
		RECT	15.575 26.575 15.625 26.705 ;
		RECT	15.575 24.155 15.625 24.285 ;
		RECT	20.495 26.575 20.545 26.705 ;
		RECT	20.495 24.155 20.545 24.285 ;
		RECT	15.775 26.575 15.825 26.705 ;
		RECT	15.775 24.155 15.825 24.285 ;
		RECT	20.295 26.575 20.345 26.705 ;
		RECT	20.295 24.155 20.345 24.285 ;
		RECT	15.375 23.465 15.425 23.595 ;
		RECT	20.695 23.465 20.745 23.595 ;
		RECT	15.575 23.695 15.625 23.825 ;
		RECT	15.575 21.275 15.625 21.405 ;
		RECT	20.495 23.695 20.545 23.825 ;
		RECT	20.495 21.275 20.545 21.405 ;
		RECT	15.775 23.695 15.825 23.825 ;
		RECT	15.775 21.275 15.825 21.405 ;
		RECT	20.295 23.695 20.345 23.825 ;
		RECT	20.295 21.275 20.345 21.405 ;
		RECT	15.375 20.585 15.425 20.715 ;
		RECT	20.695 20.585 20.745 20.715 ;
		RECT	15.575 20.815 15.625 20.945 ;
		RECT	15.575 18.395 15.625 18.525 ;
		RECT	20.495 20.815 20.545 20.945 ;
		RECT	20.495 18.395 20.545 18.525 ;
		RECT	15.775 20.815 15.825 20.945 ;
		RECT	15.775 18.395 15.825 18.525 ;
		RECT	20.295 20.815 20.345 20.945 ;
		RECT	20.295 18.395 20.345 18.525 ;
		RECT	15.375 17.705 15.425 17.835 ;
		RECT	20.695 17.705 20.745 17.835 ;
		RECT	15.575 17.935 15.625 18.065 ;
		RECT	15.575 15.515 15.625 15.645 ;
		RECT	20.495 17.935 20.545 18.065 ;
		RECT	20.495 15.515 20.545 15.645 ;
		RECT	15.775 17.935 15.825 18.065 ;
		RECT	15.775 15.515 15.825 15.645 ;
		RECT	20.295 17.935 20.345 18.065 ;
		RECT	20.295 15.515 20.345 15.645 ;
		RECT	15.375 14.825 15.425 14.955 ;
		RECT	20.695 14.825 20.745 14.955 ;
		RECT	15.575 15.055 15.625 15.185 ;
		RECT	15.575 12.635 15.625 12.765 ;
		RECT	20.495 15.055 20.545 15.185 ;
		RECT	20.495 12.635 20.545 12.765 ;
		RECT	15.775 15.055 15.825 15.185 ;
		RECT	15.775 12.635 15.825 12.765 ;
		RECT	20.295 15.055 20.345 15.185 ;
		RECT	20.295 12.635 20.345 12.765 ;
		RECT	15.375 167.465 15.425 167.595 ;
		RECT	20.695 167.465 20.745 167.595 ;
		RECT	15.575 167.695 15.625 167.825 ;
		RECT	15.575 165.275 15.625 165.405 ;
		RECT	20.495 167.695 20.545 167.825 ;
		RECT	20.495 165.275 20.545 165.405 ;
		RECT	15.775 167.695 15.825 167.825 ;
		RECT	15.775 165.275 15.825 165.405 ;
		RECT	20.295 167.695 20.345 167.825 ;
		RECT	20.295 165.275 20.345 165.405 ;
		RECT	15.375 11.945 15.425 12.075 ;
		RECT	20.695 11.945 20.745 12.075 ;
		RECT	15.575 12.175 15.625 12.305 ;
		RECT	15.575 9.755 15.625 9.885 ;
		RECT	20.495 12.175 20.545 12.305 ;
		RECT	20.495 9.755 20.545 9.885 ;
		RECT	15.775 12.175 15.825 12.305 ;
		RECT	15.775 9.755 15.825 9.885 ;
		RECT	20.295 12.175 20.345 12.305 ;
		RECT	20.295 9.755 20.345 9.885 ;
		RECT	15.375 9.065 15.425 9.195 ;
		RECT	20.695 9.065 20.745 9.195 ;
		RECT	15.575 9.295 15.625 9.425 ;
		RECT	15.575 6.875 15.625 7.005 ;
		RECT	20.495 9.295 20.545 9.425 ;
		RECT	20.495 6.875 20.545 7.005 ;
		RECT	15.775 9.295 15.825 9.425 ;
		RECT	15.775 6.875 15.825 7.005 ;
		RECT	20.295 9.295 20.345 9.425 ;
		RECT	20.295 6.875 20.345 7.005 ;
		RECT	15.375 6.185 15.425 6.315 ;
		RECT	20.695 6.185 20.745 6.315 ;
		RECT	15.575 6.415 15.625 6.545 ;
		RECT	15.575 3.995 15.625 4.125 ;
		RECT	20.495 6.415 20.545 6.545 ;
		RECT	20.495 3.995 20.545 4.125 ;
		RECT	15.775 6.415 15.825 6.545 ;
		RECT	15.775 3.995 15.825 4.125 ;
		RECT	20.295 6.415 20.345 6.545 ;
		RECT	20.295 3.995 20.345 4.125 ;
		RECT	15.375 164.585 15.425 164.715 ;
		RECT	20.695 164.585 20.745 164.715 ;
		RECT	15.575 164.815 15.625 164.945 ;
		RECT	15.575 162.395 15.625 162.525 ;
		RECT	20.495 164.815 20.545 164.945 ;
		RECT	20.495 162.395 20.545 162.525 ;
		RECT	15.775 164.815 15.825 164.945 ;
		RECT	15.775 162.395 15.825 162.525 ;
		RECT	20.295 164.815 20.345 164.945 ;
		RECT	20.295 162.395 20.345 162.525 ;
		RECT	15.375 161.705 15.425 161.835 ;
		RECT	20.695 161.705 20.745 161.835 ;
		RECT	15.575 161.935 15.625 162.065 ;
		RECT	15.575 159.515 15.625 159.645 ;
		RECT	20.495 161.935 20.545 162.065 ;
		RECT	20.495 159.515 20.545 159.645 ;
		RECT	15.775 161.935 15.825 162.065 ;
		RECT	15.775 159.515 15.825 159.645 ;
		RECT	20.295 161.935 20.345 162.065 ;
		RECT	20.295 159.515 20.345 159.645 ;
		RECT	15.375 158.825 15.425 158.955 ;
		RECT	20.695 158.825 20.745 158.955 ;
		RECT	15.575 159.055 15.625 159.185 ;
		RECT	15.575 156.635 15.625 156.765 ;
		RECT	20.495 159.055 20.545 159.185 ;
		RECT	20.495 156.635 20.545 156.765 ;
		RECT	15.775 159.055 15.825 159.185 ;
		RECT	15.775 156.635 15.825 156.765 ;
		RECT	20.295 159.055 20.345 159.185 ;
		RECT	20.295 156.635 20.345 156.765 ;
		RECT	21.025 182.095 21.075 182.225 ;
		RECT	20.895 182.095 20.945 182.225 ;
		RECT	21.815 181.865 21.865 181.995 ;
		RECT	21.685 181.865 21.735 181.995 ;
		RECT	21.025 179.675 21.075 179.805 ;
		RECT	20.895 179.675 20.945 179.805 ;
		RECT	21.24 179.445 21.29 179.575 ;
		RECT	21.025 156.175 21.075 156.305 ;
		RECT	20.895 156.175 20.945 156.305 ;
		RECT	21.815 155.945 21.865 156.075 ;
		RECT	21.685 155.945 21.735 156.075 ;
		RECT	21.025 153.755 21.075 153.885 ;
		RECT	20.895 153.755 20.945 153.885 ;
		RECT	21.24 153.525 21.29 153.655 ;
		RECT	21.025 153.295 21.075 153.425 ;
		RECT	20.895 153.295 20.945 153.425 ;
		RECT	21.815 153.065 21.865 153.195 ;
		RECT	21.685 153.065 21.735 153.195 ;
		RECT	21.025 150.875 21.075 151.005 ;
		RECT	20.895 150.875 20.945 151.005 ;
		RECT	21.24 150.645 21.29 150.775 ;
		RECT	21.025 150.415 21.075 150.545 ;
		RECT	20.895 150.415 20.945 150.545 ;
		RECT	21.815 150.185 21.865 150.315 ;
		RECT	21.685 150.185 21.735 150.315 ;
		RECT	21.025 147.995 21.075 148.125 ;
		RECT	20.895 147.995 20.945 148.125 ;
		RECT	21.24 147.765 21.29 147.895 ;
		RECT	21.025 147.535 21.075 147.665 ;
		RECT	20.895 147.535 20.945 147.665 ;
		RECT	21.815 147.305 21.865 147.435 ;
		RECT	21.685 147.305 21.735 147.435 ;
		RECT	21.025 145.115 21.075 145.245 ;
		RECT	20.895 145.115 20.945 145.245 ;
		RECT	21.24 144.885 21.29 145.015 ;
		RECT	21.025 144.655 21.075 144.785 ;
		RECT	20.895 144.655 20.945 144.785 ;
		RECT	21.815 144.425 21.865 144.555 ;
		RECT	21.685 144.425 21.735 144.555 ;
		RECT	21.025 142.235 21.075 142.365 ;
		RECT	20.895 142.235 20.945 142.365 ;
		RECT	21.24 142.005 21.29 142.135 ;
		RECT	21.025 141.775 21.075 141.905 ;
		RECT	20.895 141.775 20.945 141.905 ;
		RECT	21.815 141.545 21.865 141.675 ;
		RECT	21.685 141.545 21.735 141.675 ;
		RECT	21.025 139.355 21.075 139.485 ;
		RECT	20.895 139.355 20.945 139.485 ;
		RECT	21.24 139.125 21.29 139.255 ;
		RECT	21.025 138.895 21.075 139.025 ;
		RECT	20.895 138.895 20.945 139.025 ;
		RECT	21.815 138.665 21.865 138.795 ;
		RECT	21.685 138.665 21.735 138.795 ;
		RECT	21.025 136.475 21.075 136.605 ;
		RECT	20.895 136.475 20.945 136.605 ;
		RECT	21.24 136.245 21.29 136.375 ;
		RECT	21.025 136.015 21.075 136.145 ;
		RECT	20.895 136.015 20.945 136.145 ;
		RECT	21.815 135.785 21.865 135.915 ;
		RECT	21.685 135.785 21.735 135.915 ;
		RECT	21.025 133.595 21.075 133.725 ;
		RECT	20.895 133.595 20.945 133.725 ;
		RECT	21.24 133.365 21.29 133.495 ;
		RECT	21.025 133.135 21.075 133.265 ;
		RECT	20.895 133.135 20.945 133.265 ;
		RECT	21.815 132.905 21.865 133.035 ;
		RECT	21.685 132.905 21.735 133.035 ;
		RECT	21.025 130.715 21.075 130.845 ;
		RECT	20.895 130.715 20.945 130.845 ;
		RECT	21.24 130.485 21.29 130.615 ;
		RECT	21.025 130.255 21.075 130.385 ;
		RECT	20.895 130.255 20.945 130.385 ;
		RECT	21.815 130.025 21.865 130.155 ;
		RECT	21.685 130.025 21.735 130.155 ;
		RECT	21.025 127.835 21.075 127.965 ;
		RECT	20.895 127.835 20.945 127.965 ;
		RECT	21.24 127.605 21.29 127.735 ;
		RECT	21.025 179.215 21.075 179.345 ;
		RECT	20.895 179.215 20.945 179.345 ;
		RECT	21.815 178.985 21.865 179.115 ;
		RECT	21.685 178.985 21.735 179.115 ;
		RECT	21.025 176.795 21.075 176.925 ;
		RECT	20.895 176.795 20.945 176.925 ;
		RECT	21.24 176.565 21.29 176.695 ;
		RECT	21.025 127.375 21.075 127.505 ;
		RECT	20.895 127.375 20.945 127.505 ;
		RECT	21.815 127.145 21.865 127.275 ;
		RECT	21.685 127.145 21.735 127.275 ;
		RECT	21.025 124.955 21.075 125.085 ;
		RECT	20.895 124.955 20.945 125.085 ;
		RECT	21.24 124.725 21.29 124.855 ;
		RECT	21.025 124.495 21.075 124.625 ;
		RECT	20.895 124.495 20.945 124.625 ;
		RECT	21.815 124.265 21.865 124.395 ;
		RECT	21.685 124.265 21.735 124.395 ;
		RECT	21.025 122.075 21.075 122.205 ;
		RECT	20.895 122.075 20.945 122.205 ;
		RECT	21.24 121.845 21.29 121.975 ;
		RECT	21.025 121.615 21.075 121.745 ;
		RECT	20.895 121.615 20.945 121.745 ;
		RECT	21.815 121.385 21.865 121.515 ;
		RECT	21.685 121.385 21.735 121.515 ;
		RECT	21.025 119.195 21.075 119.325 ;
		RECT	20.895 119.195 20.945 119.325 ;
		RECT	21.24 118.965 21.29 119.095 ;
		RECT	21.025 118.735 21.075 118.865 ;
		RECT	20.895 118.735 20.945 118.865 ;
		RECT	21.815 118.505 21.865 118.635 ;
		RECT	21.685 118.505 21.735 118.635 ;
		RECT	21.025 116.315 21.075 116.445 ;
		RECT	20.895 116.315 20.945 116.445 ;
		RECT	21.24 116.085 21.29 116.215 ;
		RECT	21.025 115.855 21.075 115.985 ;
		RECT	20.895 115.855 20.945 115.985 ;
		RECT	21.815 115.625 21.865 115.755 ;
		RECT	21.685 115.625 21.735 115.755 ;
		RECT	21.025 113.435 21.075 113.565 ;
		RECT	20.895 113.435 20.945 113.565 ;
		RECT	21.24 113.205 21.29 113.335 ;
		RECT	21.025 112.975 21.075 113.105 ;
		RECT	20.895 112.975 20.945 113.105 ;
		RECT	21.815 112.745 21.865 112.875 ;
		RECT	21.685 112.745 21.735 112.875 ;
		RECT	21.025 110.555 21.075 110.685 ;
		RECT	20.895 110.555 20.945 110.685 ;
		RECT	21.24 110.325 21.29 110.455 ;
		RECT	21.025 110.095 21.075 110.225 ;
		RECT	20.895 110.095 20.945 110.225 ;
		RECT	21.815 109.865 21.865 109.995 ;
		RECT	21.685 109.865 21.735 109.995 ;
		RECT	21.025 107.675 21.075 107.805 ;
		RECT	20.895 107.675 20.945 107.805 ;
		RECT	21.24 107.445 21.29 107.575 ;
		RECT	21.025 107.215 21.075 107.345 ;
		RECT	20.895 107.215 20.945 107.345 ;
		RECT	21.815 106.985 21.865 107.115 ;
		RECT	21.685 106.985 21.735 107.115 ;
		RECT	21.025 104.795 21.075 104.925 ;
		RECT	20.895 104.795 20.945 104.925 ;
		RECT	21.24 104.565 21.29 104.695 ;
		RECT	21.025 104.335 21.075 104.465 ;
		RECT	20.895 104.335 20.945 104.465 ;
		RECT	21.815 104.105 21.865 104.235 ;
		RECT	21.685 104.105 21.735 104.235 ;
		RECT	21.025 101.915 21.075 102.045 ;
		RECT	20.895 101.915 20.945 102.045 ;
		RECT	21.24 101.685 21.29 101.815 ;
		RECT	21.025 101.455 21.075 101.585 ;
		RECT	20.895 101.455 20.945 101.585 ;
		RECT	21.815 101.225 21.865 101.355 ;
		RECT	21.685 101.225 21.735 101.355 ;
		RECT	21.025 99.035 21.075 99.165 ;
		RECT	20.895 99.035 20.945 99.165 ;
		RECT	21.24 98.805 21.29 98.935 ;
		RECT	21.025 176.335 21.075 176.465 ;
		RECT	20.895 176.335 20.945 176.465 ;
		RECT	21.815 176.105 21.865 176.235 ;
		RECT	21.685 176.105 21.735 176.235 ;
		RECT	21.025 173.915 21.075 174.045 ;
		RECT	20.895 173.915 20.945 174.045 ;
		RECT	21.24 173.685 21.29 173.815 ;
		RECT	21.025 98.575 21.075 98.705 ;
		RECT	20.895 98.575 20.945 98.705 ;
		RECT	21.815 98.345 21.865 98.475 ;
		RECT	21.685 98.345 21.735 98.475 ;
		RECT	21.025 96.155 21.075 96.285 ;
		RECT	20.895 96.155 20.945 96.285 ;
		RECT	21.24 95.925 21.29 96.055 ;
		RECT	21.025 95.695 21.075 95.825 ;
		RECT	20.895 95.695 20.945 95.825 ;
		RECT	21.815 95.465 21.865 95.595 ;
		RECT	21.685 95.465 21.735 95.595 ;
		RECT	21.025 93.275 21.075 93.405 ;
		RECT	20.895 93.275 20.945 93.405 ;
		RECT	21.24 93.045 21.29 93.175 ;
		RECT	21.025 92.815 21.075 92.945 ;
		RECT	20.895 92.815 20.945 92.945 ;
		RECT	21.815 92.585 21.865 92.715 ;
		RECT	21.685 92.585 21.735 92.715 ;
		RECT	21.025 90.395 21.075 90.525 ;
		RECT	20.895 90.395 20.945 90.525 ;
		RECT	21.24 90.165 21.29 90.295 ;
		RECT	21.025 89.935 21.075 90.065 ;
		RECT	20.895 89.935 20.945 90.065 ;
		RECT	21.815 89.705 21.865 89.835 ;
		RECT	21.685 89.705 21.735 89.835 ;
		RECT	21.025 87.515 21.075 87.645 ;
		RECT	20.895 87.515 20.945 87.645 ;
		RECT	21.24 87.285 21.29 87.415 ;
		RECT	21.025 87.055 21.075 87.185 ;
		RECT	20.895 87.055 20.945 87.185 ;
		RECT	21.815 86.825 21.865 86.955 ;
		RECT	21.685 86.825 21.735 86.955 ;
		RECT	21.025 84.635 21.075 84.765 ;
		RECT	20.895 84.635 20.945 84.765 ;
		RECT	21.24 84.405 21.29 84.535 ;
		RECT	21.025 84.175 21.075 84.305 ;
		RECT	20.895 84.175 20.945 84.305 ;
		RECT	21.815 83.945 21.865 84.075 ;
		RECT	21.685 83.945 21.735 84.075 ;
		RECT	21.025 81.755 21.075 81.885 ;
		RECT	20.895 81.755 20.945 81.885 ;
		RECT	21.24 81.525 21.29 81.655 ;
		RECT	21.025 81.295 21.075 81.425 ;
		RECT	20.895 81.295 20.945 81.425 ;
		RECT	21.815 81.065 21.865 81.195 ;
		RECT	21.685 81.065 21.735 81.195 ;
		RECT	21.025 78.875 21.075 79.005 ;
		RECT	20.895 78.875 20.945 79.005 ;
		RECT	21.24 78.645 21.29 78.775 ;
		RECT	21.025 78.415 21.075 78.545 ;
		RECT	20.895 78.415 20.945 78.545 ;
		RECT	21.815 78.185 21.865 78.315 ;
		RECT	21.685 78.185 21.735 78.315 ;
		RECT	21.025 75.995 21.075 76.125 ;
		RECT	20.895 75.995 20.945 76.125 ;
		RECT	21.24 75.765 21.29 75.895 ;
		RECT	21.025 75.535 21.075 75.665 ;
		RECT	20.895 75.535 20.945 75.665 ;
		RECT	21.815 75.305 21.865 75.435 ;
		RECT	21.685 75.305 21.735 75.435 ;
		RECT	21.025 73.115 21.075 73.245 ;
		RECT	20.895 73.115 20.945 73.245 ;
		RECT	21.24 72.885 21.29 73.015 ;
		RECT	21.025 72.655 21.075 72.785 ;
		RECT	20.895 72.655 20.945 72.785 ;
		RECT	21.815 72.425 21.865 72.555 ;
		RECT	21.685 72.425 21.735 72.555 ;
		RECT	21.025 70.235 21.075 70.365 ;
		RECT	20.895 70.235 20.945 70.365 ;
		RECT	21.24 70.005 21.29 70.135 ;
		RECT	21.025 173.455 21.075 173.585 ;
		RECT	20.895 173.455 20.945 173.585 ;
		RECT	21.815 173.225 21.865 173.355 ;
		RECT	21.685 173.225 21.735 173.355 ;
		RECT	21.025 171.035 21.075 171.165 ;
		RECT	20.895 171.035 20.945 171.165 ;
		RECT	21.24 170.805 21.29 170.935 ;
		RECT	21.025 69.775 21.075 69.905 ;
		RECT	20.895 69.775 20.945 69.905 ;
		RECT	21.815 69.545 21.865 69.675 ;
		RECT	21.685 69.545 21.735 69.675 ;
		RECT	21.025 67.355 21.075 67.485 ;
		RECT	20.895 67.355 20.945 67.485 ;
		RECT	21.24 67.125 21.29 67.255 ;
		RECT	21.025 66.895 21.075 67.025 ;
		RECT	20.895 66.895 20.945 67.025 ;
		RECT	21.815 66.665 21.865 66.795 ;
		RECT	21.685 66.665 21.735 66.795 ;
		RECT	21.025 64.475 21.075 64.605 ;
		RECT	20.895 64.475 20.945 64.605 ;
		RECT	21.24 64.245 21.29 64.375 ;
		RECT	21.025 64.015 21.075 64.145 ;
		RECT	20.895 64.015 20.945 64.145 ;
		RECT	21.815 63.785 21.865 63.915 ;
		RECT	21.685 63.785 21.735 63.915 ;
		RECT	21.025 61.595 21.075 61.725 ;
		RECT	20.895 61.595 20.945 61.725 ;
		RECT	21.24 61.365 21.29 61.495 ;
		RECT	21.025 61.135 21.075 61.265 ;
		RECT	20.895 61.135 20.945 61.265 ;
		RECT	21.815 60.905 21.865 61.035 ;
		RECT	21.685 60.905 21.735 61.035 ;
		RECT	21.025 58.715 21.075 58.845 ;
		RECT	20.895 58.715 20.945 58.845 ;
		RECT	21.24 58.485 21.29 58.615 ;
		RECT	21.025 58.255 21.075 58.385 ;
		RECT	20.895 58.255 20.945 58.385 ;
		RECT	21.815 58.025 21.865 58.155 ;
		RECT	21.685 58.025 21.735 58.155 ;
		RECT	21.025 55.835 21.075 55.965 ;
		RECT	20.895 55.835 20.945 55.965 ;
		RECT	21.24 55.605 21.29 55.735 ;
		RECT	21.025 55.375 21.075 55.505 ;
		RECT	20.895 55.375 20.945 55.505 ;
		RECT	21.815 55.145 21.865 55.275 ;
		RECT	21.685 55.145 21.735 55.275 ;
		RECT	21.025 52.955 21.075 53.085 ;
		RECT	20.895 52.955 20.945 53.085 ;
		RECT	21.24 52.725 21.29 52.855 ;
		RECT	21.025 52.495 21.075 52.625 ;
		RECT	20.895 52.495 20.945 52.625 ;
		RECT	21.815 52.265 21.865 52.395 ;
		RECT	21.685 52.265 21.735 52.395 ;
		RECT	21.025 50.075 21.075 50.205 ;
		RECT	20.895 50.075 20.945 50.205 ;
		RECT	21.24 49.845 21.29 49.975 ;
		RECT	21.025 49.615 21.075 49.745 ;
		RECT	20.895 49.615 20.945 49.745 ;
		RECT	21.815 49.385 21.865 49.515 ;
		RECT	21.685 49.385 21.735 49.515 ;
		RECT	21.025 47.195 21.075 47.325 ;
		RECT	20.895 47.195 20.945 47.325 ;
		RECT	21.24 46.965 21.29 47.095 ;
		RECT	21.025 46.735 21.075 46.865 ;
		RECT	20.895 46.735 20.945 46.865 ;
		RECT	21.815 46.505 21.865 46.635 ;
		RECT	21.685 46.505 21.735 46.635 ;
		RECT	21.025 44.315 21.075 44.445 ;
		RECT	20.895 44.315 20.945 44.445 ;
		RECT	21.24 44.085 21.29 44.215 ;
		RECT	21.025 43.855 21.075 43.985 ;
		RECT	20.895 43.855 20.945 43.985 ;
		RECT	21.815 43.625 21.865 43.755 ;
		RECT	21.685 43.625 21.735 43.755 ;
		RECT	21.025 41.435 21.075 41.565 ;
		RECT	20.895 41.435 20.945 41.565 ;
		RECT	21.24 41.205 21.29 41.335 ;
		RECT	21.025 170.575 21.075 170.705 ;
		RECT	20.895 170.575 20.945 170.705 ;
		RECT	21.815 170.345 21.865 170.475 ;
		RECT	21.685 170.345 21.735 170.475 ;
		RECT	21.025 168.155 21.075 168.285 ;
		RECT	20.895 168.155 20.945 168.285 ;
		RECT	21.24 167.925 21.29 168.055 ;
		RECT	21.025 40.975 21.075 41.105 ;
		RECT	20.895 40.975 20.945 41.105 ;
		RECT	21.815 40.745 21.865 40.875 ;
		RECT	21.685 40.745 21.735 40.875 ;
		RECT	21.025 38.555 21.075 38.685 ;
		RECT	20.895 38.555 20.945 38.685 ;
		RECT	21.24 38.325 21.29 38.455 ;
		RECT	21.025 38.095 21.075 38.225 ;
		RECT	20.895 38.095 20.945 38.225 ;
		RECT	21.815 37.865 21.865 37.995 ;
		RECT	21.685 37.865 21.735 37.995 ;
		RECT	21.025 35.675 21.075 35.805 ;
		RECT	20.895 35.675 20.945 35.805 ;
		RECT	21.24 35.445 21.29 35.575 ;
		RECT	21.025 35.215 21.075 35.345 ;
		RECT	20.895 35.215 20.945 35.345 ;
		RECT	21.815 34.985 21.865 35.115 ;
		RECT	21.685 34.985 21.735 35.115 ;
		RECT	21.025 32.795 21.075 32.925 ;
		RECT	20.895 32.795 20.945 32.925 ;
		RECT	21.24 32.565 21.29 32.695 ;
		RECT	21.025 32.335 21.075 32.465 ;
		RECT	20.895 32.335 20.945 32.465 ;
		RECT	21.815 32.105 21.865 32.235 ;
		RECT	21.685 32.105 21.735 32.235 ;
		RECT	21.025 29.915 21.075 30.045 ;
		RECT	20.895 29.915 20.945 30.045 ;
		RECT	21.24 29.685 21.29 29.815 ;
		RECT	21.025 29.455 21.075 29.585 ;
		RECT	20.895 29.455 20.945 29.585 ;
		RECT	21.815 29.225 21.865 29.355 ;
		RECT	21.685 29.225 21.735 29.355 ;
		RECT	21.025 27.035 21.075 27.165 ;
		RECT	20.895 27.035 20.945 27.165 ;
		RECT	21.24 26.805 21.29 26.935 ;
		RECT	21.025 26.575 21.075 26.705 ;
		RECT	20.895 26.575 20.945 26.705 ;
		RECT	21.815 26.345 21.865 26.475 ;
		RECT	21.685 26.345 21.735 26.475 ;
		RECT	21.025 24.155 21.075 24.285 ;
		RECT	20.895 24.155 20.945 24.285 ;
		RECT	21.24 23.925 21.29 24.055 ;
		RECT	21.025 23.695 21.075 23.825 ;
		RECT	20.895 23.695 20.945 23.825 ;
		RECT	21.815 23.465 21.865 23.595 ;
		RECT	21.685 23.465 21.735 23.595 ;
		RECT	21.025 21.275 21.075 21.405 ;
		RECT	20.895 21.275 20.945 21.405 ;
		RECT	21.24 21.045 21.29 21.175 ;
		RECT	21.025 20.815 21.075 20.945 ;
		RECT	20.895 20.815 20.945 20.945 ;
		RECT	21.815 20.585 21.865 20.715 ;
		RECT	21.685 20.585 21.735 20.715 ;
		RECT	21.025 18.395 21.075 18.525 ;
		RECT	20.895 18.395 20.945 18.525 ;
		RECT	21.24 18.165 21.29 18.295 ;
		RECT	21.025 17.935 21.075 18.065 ;
		RECT	20.895 17.935 20.945 18.065 ;
		RECT	21.815 17.705 21.865 17.835 ;
		RECT	21.685 17.705 21.735 17.835 ;
		RECT	21.025 15.515 21.075 15.645 ;
		RECT	20.895 15.515 20.945 15.645 ;
		RECT	21.24 15.285 21.29 15.415 ;
		RECT	21.025 15.055 21.075 15.185 ;
		RECT	20.895 15.055 20.945 15.185 ;
		RECT	21.815 14.825 21.865 14.955 ;
		RECT	21.685 14.825 21.735 14.955 ;
		RECT	21.025 12.635 21.075 12.765 ;
		RECT	20.895 12.635 20.945 12.765 ;
		RECT	21.24 12.405 21.29 12.535 ;
		RECT	21.025 167.695 21.075 167.825 ;
		RECT	20.895 167.695 20.945 167.825 ;
		RECT	21.815 167.465 21.865 167.595 ;
		RECT	21.685 167.465 21.735 167.595 ;
		RECT	21.025 165.275 21.075 165.405 ;
		RECT	20.895 165.275 20.945 165.405 ;
		RECT	21.24 165.045 21.29 165.175 ;
		RECT	21.025 12.175 21.075 12.305 ;
		RECT	20.895 12.175 20.945 12.305 ;
		RECT	21.815 11.945 21.865 12.075 ;
		RECT	21.685 11.945 21.735 12.075 ;
		RECT	21.025 9.755 21.075 9.885 ;
		RECT	20.895 9.755 20.945 9.885 ;
		RECT	21.24 9.525 21.29 9.655 ;
		RECT	21.025 9.295 21.075 9.425 ;
		RECT	20.895 9.295 20.945 9.425 ;
		RECT	21.815 9.065 21.865 9.195 ;
		RECT	21.685 9.065 21.735 9.195 ;
		RECT	21.025 6.875 21.075 7.005 ;
		RECT	20.895 6.875 20.945 7.005 ;
		RECT	21.24 6.645 21.29 6.775 ;
		RECT	21.025 6.415 21.075 6.545 ;
		RECT	20.895 6.415 20.945 6.545 ;
		RECT	21.815 6.185 21.865 6.315 ;
		RECT	21.685 6.185 21.735 6.315 ;
		RECT	21.025 3.995 21.075 4.125 ;
		RECT	20.895 3.995 20.945 4.125 ;
		RECT	21.24 3.765 21.29 3.895 ;
		RECT	21.025 164.815 21.075 164.945 ;
		RECT	20.895 164.815 20.945 164.945 ;
		RECT	21.815 164.585 21.865 164.715 ;
		RECT	21.685 164.585 21.735 164.715 ;
		RECT	21.025 162.395 21.075 162.525 ;
		RECT	20.895 162.395 20.945 162.525 ;
		RECT	21.24 162.165 21.29 162.295 ;
		RECT	21.025 161.935 21.075 162.065 ;
		RECT	20.895 161.935 20.945 162.065 ;
		RECT	21.815 161.705 21.865 161.835 ;
		RECT	21.685 161.705 21.735 161.835 ;
		RECT	21.025 159.515 21.075 159.645 ;
		RECT	20.895 159.515 20.945 159.645 ;
		RECT	21.24 159.285 21.29 159.415 ;
		RECT	21.025 159.055 21.075 159.185 ;
		RECT	20.895 159.055 20.945 159.185 ;
		RECT	21.815 158.825 21.865 158.955 ;
		RECT	21.685 158.825 21.735 158.955 ;
		RECT	21.025 156.635 21.075 156.765 ;
		RECT	20.895 156.635 20.945 156.765 ;
		RECT	21.24 156.405 21.29 156.535 ;
		RECT	21.025 3.535 21.075 3.665 ;
		RECT	20.895 3.535 20.945 3.665 ;
		RECT	21.815 3.305 21.865 3.435 ;
		RECT	21.685 3.305 21.735 3.435 ;
		RECT	21.025 1.115 21.075 1.245 ;
		RECT	20.895 1.115 20.945 1.245 ;
		RECT	21.24 0.885 21.29 1.015 ;
		RECT	21.025 184.975 21.075 185.105 ;
		RECT	20.895 184.975 20.945 185.105 ;
		RECT	21.815 184.745 21.865 184.875 ;
		RECT	21.685 184.745 21.735 184.875 ;
		RECT	21.025 182.555 21.075 182.685 ;
		RECT	20.895 182.555 20.945 182.685 ;
		RECT	21.24 182.325 21.29 182.455 ;
		RECT	15.375 411.425 15.425 411.555 ;
		RECT	20.695 411.425 20.745 411.555 ;
		RECT	15.575 411.195 15.625 411.325 ;
		RECT	15.575 413.615 15.625 413.745 ;
		RECT	20.495 411.195 20.545 411.325 ;
		RECT	20.495 413.615 20.545 413.745 ;
		RECT	15.775 411.195 15.825 411.325 ;
		RECT	15.775 413.615 15.825 413.745 ;
		RECT	20.295 411.195 20.345 411.325 ;
		RECT	20.295 413.615 20.345 413.745 ;
		RECT	15.375 229.985 15.425 230.115 ;
		RECT	20.695 229.985 20.745 230.115 ;
		RECT	15.575 229.755 15.625 229.885 ;
		RECT	15.575 232.175 15.625 232.305 ;
		RECT	20.495 229.755 20.545 229.885 ;
		RECT	20.495 232.175 20.545 232.305 ;
		RECT	15.775 229.755 15.825 229.885 ;
		RECT	15.775 232.175 15.825 232.305 ;
		RECT	20.295 229.755 20.345 229.885 ;
		RECT	20.295 232.175 20.345 232.305 ;
		RECT	15.375 232.865 15.425 232.995 ;
		RECT	20.695 232.865 20.745 232.995 ;
		RECT	15.575 232.635 15.625 232.765 ;
		RECT	15.575 235.055 15.625 235.185 ;
		RECT	20.495 232.635 20.545 232.765 ;
		RECT	20.495 235.055 20.545 235.185 ;
		RECT	15.775 232.635 15.825 232.765 ;
		RECT	15.775 235.055 15.825 235.185 ;
		RECT	20.295 232.635 20.345 232.765 ;
		RECT	20.295 235.055 20.345 235.185 ;
		RECT	15.375 258.785 15.425 258.915 ;
		RECT	20.695 258.785 20.745 258.915 ;
		RECT	15.575 258.555 15.625 258.685 ;
		RECT	15.575 260.975 15.625 261.105 ;
		RECT	20.495 258.555 20.545 258.685 ;
		RECT	20.495 260.975 20.545 261.105 ;
		RECT	15.775 258.555 15.825 258.685 ;
		RECT	15.775 260.975 15.825 261.105 ;
		RECT	20.295 258.555 20.345 258.685 ;
		RECT	20.295 260.975 20.345 261.105 ;
		RECT	15.375 261.665 15.425 261.795 ;
		RECT	20.695 261.665 20.745 261.795 ;
		RECT	15.575 261.435 15.625 261.565 ;
		RECT	15.575 263.855 15.625 263.985 ;
		RECT	20.495 261.435 20.545 261.565 ;
		RECT	20.495 263.855 20.545 263.985 ;
		RECT	15.775 261.435 15.825 261.565 ;
		RECT	15.775 263.855 15.825 263.985 ;
		RECT	20.295 261.435 20.345 261.565 ;
		RECT	20.295 263.855 20.345 263.985 ;
		RECT	15.375 264.545 15.425 264.675 ;
		RECT	20.695 264.545 20.745 264.675 ;
		RECT	15.575 264.315 15.625 264.445 ;
		RECT	15.575 266.735 15.625 266.865 ;
		RECT	20.495 264.315 20.545 264.445 ;
		RECT	20.495 266.735 20.545 266.865 ;
		RECT	15.775 264.315 15.825 264.445 ;
		RECT	15.775 266.735 15.825 266.865 ;
		RECT	20.295 264.315 20.345 264.445 ;
		RECT	20.295 266.735 20.345 266.865 ;
		RECT	15.375 267.425 15.425 267.555 ;
		RECT	20.695 267.425 20.745 267.555 ;
		RECT	15.575 267.195 15.625 267.325 ;
		RECT	15.575 269.615 15.625 269.745 ;
		RECT	20.495 267.195 20.545 267.325 ;
		RECT	20.495 269.615 20.545 269.745 ;
		RECT	15.775 267.195 15.825 267.325 ;
		RECT	15.775 269.615 15.825 269.745 ;
		RECT	20.295 267.195 20.345 267.325 ;
		RECT	20.295 269.615 20.345 269.745 ;
		RECT	15.375 270.305 15.425 270.435 ;
		RECT	20.695 270.305 20.745 270.435 ;
		RECT	15.575 270.075 15.625 270.205 ;
		RECT	15.575 272.495 15.625 272.625 ;
		RECT	20.495 270.075 20.545 270.205 ;
		RECT	20.495 272.495 20.545 272.625 ;
		RECT	15.775 270.075 15.825 270.205 ;
		RECT	15.775 272.495 15.825 272.625 ;
		RECT	20.295 270.075 20.345 270.205 ;
		RECT	20.295 272.495 20.345 272.625 ;
		RECT	15.375 273.185 15.425 273.315 ;
		RECT	20.695 273.185 20.745 273.315 ;
		RECT	15.575 272.955 15.625 273.085 ;
		RECT	15.575 275.375 15.625 275.505 ;
		RECT	20.495 272.955 20.545 273.085 ;
		RECT	20.495 275.375 20.545 275.505 ;
		RECT	15.775 272.955 15.825 273.085 ;
		RECT	15.775 275.375 15.825 275.505 ;
		RECT	20.295 272.955 20.345 273.085 ;
		RECT	20.295 275.375 20.345 275.505 ;
		RECT	15.375 276.065 15.425 276.195 ;
		RECT	20.695 276.065 20.745 276.195 ;
		RECT	15.575 275.835 15.625 275.965 ;
		RECT	15.575 278.255 15.625 278.385 ;
		RECT	20.495 275.835 20.545 275.965 ;
		RECT	20.495 278.255 20.545 278.385 ;
		RECT	15.775 275.835 15.825 275.965 ;
		RECT	15.775 278.255 15.825 278.385 ;
		RECT	20.295 275.835 20.345 275.965 ;
		RECT	20.295 278.255 20.345 278.385 ;
		RECT	15.375 278.945 15.425 279.075 ;
		RECT	20.695 278.945 20.745 279.075 ;
		RECT	15.575 278.715 15.625 278.845 ;
		RECT	15.575 281.135 15.625 281.265 ;
		RECT	20.495 278.715 20.545 278.845 ;
		RECT	20.495 281.135 20.545 281.265 ;
		RECT	15.775 278.715 15.825 278.845 ;
		RECT	15.775 281.135 15.825 281.265 ;
		RECT	20.295 278.715 20.345 278.845 ;
		RECT	20.295 281.135 20.345 281.265 ;
		RECT	15.375 281.825 15.425 281.955 ;
		RECT	20.695 281.825 20.745 281.955 ;
		RECT	15.575 281.595 15.625 281.725 ;
		RECT	15.575 284.015 15.625 284.145 ;
		RECT	20.495 281.595 20.545 281.725 ;
		RECT	20.495 284.015 20.545 284.145 ;
		RECT	15.775 281.595 15.825 281.725 ;
		RECT	15.775 284.015 15.825 284.145 ;
		RECT	20.295 281.595 20.345 281.725 ;
		RECT	20.295 284.015 20.345 284.145 ;
		RECT	15.375 284.705 15.425 284.835 ;
		RECT	20.695 284.705 20.745 284.835 ;
		RECT	15.575 284.475 15.625 284.605 ;
		RECT	15.575 286.895 15.625 287.025 ;
		RECT	20.495 284.475 20.545 284.605 ;
		RECT	20.495 286.895 20.545 287.025 ;
		RECT	15.775 284.475 15.825 284.605 ;
		RECT	15.775 286.895 15.825 287.025 ;
		RECT	20.295 284.475 20.345 284.605 ;
		RECT	20.295 286.895 20.345 287.025 ;
		RECT	15.375 235.745 15.425 235.875 ;
		RECT	20.695 235.745 20.745 235.875 ;
		RECT	15.575 235.515 15.625 235.645 ;
		RECT	15.575 237.935 15.625 238.065 ;
		RECT	20.495 235.515 20.545 235.645 ;
		RECT	20.495 237.935 20.545 238.065 ;
		RECT	15.775 235.515 15.825 235.645 ;
		RECT	15.775 237.935 15.825 238.065 ;
		RECT	20.295 235.515 20.345 235.645 ;
		RECT	20.295 237.935 20.345 238.065 ;
		RECT	15.375 287.585 15.425 287.715 ;
		RECT	20.695 287.585 20.745 287.715 ;
		RECT	15.575 287.355 15.625 287.485 ;
		RECT	15.575 289.775 15.625 289.905 ;
		RECT	20.495 287.355 20.545 287.485 ;
		RECT	20.495 289.775 20.545 289.905 ;
		RECT	15.775 287.355 15.825 287.485 ;
		RECT	15.775 289.775 15.825 289.905 ;
		RECT	20.295 287.355 20.345 287.485 ;
		RECT	20.295 289.775 20.345 289.905 ;
		RECT	15.375 290.465 15.425 290.595 ;
		RECT	20.695 290.465 20.745 290.595 ;
		RECT	15.575 290.235 15.625 290.365 ;
		RECT	15.575 292.655 15.625 292.785 ;
		RECT	20.495 290.235 20.545 290.365 ;
		RECT	20.495 292.655 20.545 292.785 ;
		RECT	15.775 290.235 15.825 290.365 ;
		RECT	15.775 292.655 15.825 292.785 ;
		RECT	20.295 290.235 20.345 290.365 ;
		RECT	20.295 292.655 20.345 292.785 ;
		RECT	15.375 293.345 15.425 293.475 ;
		RECT	20.695 293.345 20.745 293.475 ;
		RECT	15.575 293.115 15.625 293.245 ;
		RECT	15.575 295.535 15.625 295.665 ;
		RECT	20.495 293.115 20.545 293.245 ;
		RECT	20.495 295.535 20.545 295.665 ;
		RECT	15.775 293.115 15.825 293.245 ;
		RECT	15.775 295.535 15.825 295.665 ;
		RECT	20.295 293.115 20.345 293.245 ;
		RECT	20.295 295.535 20.345 295.665 ;
		RECT	15.375 296.225 15.425 296.355 ;
		RECT	20.695 296.225 20.745 296.355 ;
		RECT	15.575 295.995 15.625 296.125 ;
		RECT	15.575 298.415 15.625 298.545 ;
		RECT	20.495 295.995 20.545 296.125 ;
		RECT	20.495 298.415 20.545 298.545 ;
		RECT	15.775 295.995 15.825 296.125 ;
		RECT	15.775 298.415 15.825 298.545 ;
		RECT	20.295 295.995 20.345 296.125 ;
		RECT	20.295 298.415 20.345 298.545 ;
		RECT	15.375 299.105 15.425 299.235 ;
		RECT	20.695 299.105 20.745 299.235 ;
		RECT	15.575 298.875 15.625 299.005 ;
		RECT	15.575 301.295 15.625 301.425 ;
		RECT	20.495 298.875 20.545 299.005 ;
		RECT	20.495 301.295 20.545 301.425 ;
		RECT	15.775 298.875 15.825 299.005 ;
		RECT	15.775 301.295 15.825 301.425 ;
		RECT	20.295 298.875 20.345 299.005 ;
		RECT	20.295 301.295 20.345 301.425 ;
		RECT	15.375 301.985 15.425 302.115 ;
		RECT	20.695 301.985 20.745 302.115 ;
		RECT	15.575 301.755 15.625 301.885 ;
		RECT	15.575 304.175 15.625 304.305 ;
		RECT	20.495 301.755 20.545 301.885 ;
		RECT	20.495 304.175 20.545 304.305 ;
		RECT	15.775 301.755 15.825 301.885 ;
		RECT	15.775 304.175 15.825 304.305 ;
		RECT	20.295 301.755 20.345 301.885 ;
		RECT	20.295 304.175 20.345 304.305 ;
		RECT	15.375 304.865 15.425 304.995 ;
		RECT	20.695 304.865 20.745 304.995 ;
		RECT	15.575 304.635 15.625 304.765 ;
		RECT	15.575 307.055 15.625 307.185 ;
		RECT	20.495 304.635 20.545 304.765 ;
		RECT	20.495 307.055 20.545 307.185 ;
		RECT	15.775 304.635 15.825 304.765 ;
		RECT	15.775 307.055 15.825 307.185 ;
		RECT	20.295 304.635 20.345 304.765 ;
		RECT	20.295 307.055 20.345 307.185 ;
		RECT	15.375 307.745 15.425 307.875 ;
		RECT	20.695 307.745 20.745 307.875 ;
		RECT	15.575 307.515 15.625 307.645 ;
		RECT	15.575 309.935 15.625 310.065 ;
		RECT	20.495 307.515 20.545 307.645 ;
		RECT	20.495 309.935 20.545 310.065 ;
		RECT	15.775 307.515 15.825 307.645 ;
		RECT	15.775 309.935 15.825 310.065 ;
		RECT	20.295 307.515 20.345 307.645 ;
		RECT	20.295 309.935 20.345 310.065 ;
		RECT	15.375 310.625 15.425 310.755 ;
		RECT	20.695 310.625 20.745 310.755 ;
		RECT	15.575 310.395 15.625 310.525 ;
		RECT	15.575 312.815 15.625 312.945 ;
		RECT	20.495 310.395 20.545 310.525 ;
		RECT	20.495 312.815 20.545 312.945 ;
		RECT	15.775 310.395 15.825 310.525 ;
		RECT	15.775 312.815 15.825 312.945 ;
		RECT	20.295 310.395 20.345 310.525 ;
		RECT	20.295 312.815 20.345 312.945 ;
		RECT	15.375 313.505 15.425 313.635 ;
		RECT	20.695 313.505 20.745 313.635 ;
		RECT	15.575 313.275 15.625 313.405 ;
		RECT	15.575 315.695 15.625 315.825 ;
		RECT	20.495 313.275 20.545 313.405 ;
		RECT	20.495 315.695 20.545 315.825 ;
		RECT	15.775 313.275 15.825 313.405 ;
		RECT	15.775 315.695 15.825 315.825 ;
		RECT	20.295 313.275 20.345 313.405 ;
		RECT	20.295 315.695 20.345 315.825 ;
		RECT	15.375 238.625 15.425 238.755 ;
		RECT	20.695 238.625 20.745 238.755 ;
		RECT	15.575 238.395 15.625 238.525 ;
		RECT	15.575 240.815 15.625 240.945 ;
		RECT	20.495 238.395 20.545 238.525 ;
		RECT	20.495 240.815 20.545 240.945 ;
		RECT	15.775 238.395 15.825 238.525 ;
		RECT	15.775 240.815 15.825 240.945 ;
		RECT	20.295 238.395 20.345 238.525 ;
		RECT	20.295 240.815 20.345 240.945 ;
		RECT	15.375 316.385 15.425 316.515 ;
		RECT	20.695 316.385 20.745 316.515 ;
		RECT	15.575 316.155 15.625 316.285 ;
		RECT	15.575 318.575 15.625 318.705 ;
		RECT	20.495 316.155 20.545 316.285 ;
		RECT	20.495 318.575 20.545 318.705 ;
		RECT	15.775 316.155 15.825 316.285 ;
		RECT	15.775 318.575 15.825 318.705 ;
		RECT	20.295 316.155 20.345 316.285 ;
		RECT	20.295 318.575 20.345 318.705 ;
		RECT	15.375 319.265 15.425 319.395 ;
		RECT	20.695 319.265 20.745 319.395 ;
		RECT	15.575 319.035 15.625 319.165 ;
		RECT	15.575 321.455 15.625 321.585 ;
		RECT	20.495 319.035 20.545 319.165 ;
		RECT	20.495 321.455 20.545 321.585 ;
		RECT	15.775 319.035 15.825 319.165 ;
		RECT	15.775 321.455 15.825 321.585 ;
		RECT	20.295 319.035 20.345 319.165 ;
		RECT	20.295 321.455 20.345 321.585 ;
		RECT	15.375 322.145 15.425 322.275 ;
		RECT	20.695 322.145 20.745 322.275 ;
		RECT	15.575 321.915 15.625 322.045 ;
		RECT	15.575 324.335 15.625 324.465 ;
		RECT	20.495 321.915 20.545 322.045 ;
		RECT	20.495 324.335 20.545 324.465 ;
		RECT	15.775 321.915 15.825 322.045 ;
		RECT	15.775 324.335 15.825 324.465 ;
		RECT	20.295 321.915 20.345 322.045 ;
		RECT	20.295 324.335 20.345 324.465 ;
		RECT	15.375 325.025 15.425 325.155 ;
		RECT	20.695 325.025 20.745 325.155 ;
		RECT	15.575 324.795 15.625 324.925 ;
		RECT	15.575 327.215 15.625 327.345 ;
		RECT	20.495 324.795 20.545 324.925 ;
		RECT	20.495 327.215 20.545 327.345 ;
		RECT	15.775 324.795 15.825 324.925 ;
		RECT	15.775 327.215 15.825 327.345 ;
		RECT	20.295 324.795 20.345 324.925 ;
		RECT	20.295 327.215 20.345 327.345 ;
		RECT	15.375 327.905 15.425 328.035 ;
		RECT	20.695 327.905 20.745 328.035 ;
		RECT	15.575 327.675 15.625 327.805 ;
		RECT	15.575 330.095 15.625 330.225 ;
		RECT	20.495 327.675 20.545 327.805 ;
		RECT	20.495 330.095 20.545 330.225 ;
		RECT	15.775 327.675 15.825 327.805 ;
		RECT	15.775 330.095 15.825 330.225 ;
		RECT	20.295 327.675 20.345 327.805 ;
		RECT	20.295 330.095 20.345 330.225 ;
		RECT	15.375 330.785 15.425 330.915 ;
		RECT	20.695 330.785 20.745 330.915 ;
		RECT	15.575 330.555 15.625 330.685 ;
		RECT	15.575 332.975 15.625 333.105 ;
		RECT	20.495 330.555 20.545 330.685 ;
		RECT	20.495 332.975 20.545 333.105 ;
		RECT	15.775 330.555 15.825 330.685 ;
		RECT	15.775 332.975 15.825 333.105 ;
		RECT	20.295 330.555 20.345 330.685 ;
		RECT	20.295 332.975 20.345 333.105 ;
		RECT	15.375 333.665 15.425 333.795 ;
		RECT	20.695 333.665 20.745 333.795 ;
		RECT	15.575 333.435 15.625 333.565 ;
		RECT	15.575 335.855 15.625 335.985 ;
		RECT	20.495 333.435 20.545 333.565 ;
		RECT	20.495 335.855 20.545 335.985 ;
		RECT	15.775 333.435 15.825 333.565 ;
		RECT	15.775 335.855 15.825 335.985 ;
		RECT	20.295 333.435 20.345 333.565 ;
		RECT	20.295 335.855 20.345 335.985 ;
		RECT	15.375 336.545 15.425 336.675 ;
		RECT	20.695 336.545 20.745 336.675 ;
		RECT	15.575 336.315 15.625 336.445 ;
		RECT	15.575 338.735 15.625 338.865 ;
		RECT	20.495 336.315 20.545 336.445 ;
		RECT	20.495 338.735 20.545 338.865 ;
		RECT	15.775 336.315 15.825 336.445 ;
		RECT	15.775 338.735 15.825 338.865 ;
		RECT	20.295 336.315 20.345 336.445 ;
		RECT	20.295 338.735 20.345 338.865 ;
		RECT	15.375 339.425 15.425 339.555 ;
		RECT	20.695 339.425 20.745 339.555 ;
		RECT	15.575 339.195 15.625 339.325 ;
		RECT	15.575 341.615 15.625 341.745 ;
		RECT	20.495 339.195 20.545 339.325 ;
		RECT	20.495 341.615 20.545 341.745 ;
		RECT	15.775 339.195 15.825 339.325 ;
		RECT	15.775 341.615 15.825 341.745 ;
		RECT	20.295 339.195 20.345 339.325 ;
		RECT	20.295 341.615 20.345 341.745 ;
		RECT	15.375 342.305 15.425 342.435 ;
		RECT	20.695 342.305 20.745 342.435 ;
		RECT	15.575 342.075 15.625 342.205 ;
		RECT	15.575 344.495 15.625 344.625 ;
		RECT	20.495 342.075 20.545 342.205 ;
		RECT	20.495 344.495 20.545 344.625 ;
		RECT	15.775 342.075 15.825 342.205 ;
		RECT	15.775 344.495 15.825 344.625 ;
		RECT	20.295 342.075 20.345 342.205 ;
		RECT	20.295 344.495 20.345 344.625 ;
		RECT	15.375 241.505 15.425 241.635 ;
		RECT	20.695 241.505 20.745 241.635 ;
		RECT	15.575 241.275 15.625 241.405 ;
		RECT	15.575 243.695 15.625 243.825 ;
		RECT	20.495 241.275 20.545 241.405 ;
		RECT	20.495 243.695 20.545 243.825 ;
		RECT	15.775 241.275 15.825 241.405 ;
		RECT	15.775 243.695 15.825 243.825 ;
		RECT	20.295 241.275 20.345 241.405 ;
		RECT	20.295 243.695 20.345 243.825 ;
		RECT	15.375 345.185 15.425 345.315 ;
		RECT	20.695 345.185 20.745 345.315 ;
		RECT	15.575 344.955 15.625 345.085 ;
		RECT	15.575 347.375 15.625 347.505 ;
		RECT	20.495 344.955 20.545 345.085 ;
		RECT	20.495 347.375 20.545 347.505 ;
		RECT	15.775 344.955 15.825 345.085 ;
		RECT	15.775 347.375 15.825 347.505 ;
		RECT	20.295 344.955 20.345 345.085 ;
		RECT	20.295 347.375 20.345 347.505 ;
		RECT	15.375 348.065 15.425 348.195 ;
		RECT	20.695 348.065 20.745 348.195 ;
		RECT	15.575 347.835 15.625 347.965 ;
		RECT	15.575 350.255 15.625 350.385 ;
		RECT	20.495 347.835 20.545 347.965 ;
		RECT	20.495 350.255 20.545 350.385 ;
		RECT	15.775 347.835 15.825 347.965 ;
		RECT	15.775 350.255 15.825 350.385 ;
		RECT	20.295 347.835 20.345 347.965 ;
		RECT	20.295 350.255 20.345 350.385 ;
		RECT	15.375 350.945 15.425 351.075 ;
		RECT	20.695 350.945 20.745 351.075 ;
		RECT	15.575 350.715 15.625 350.845 ;
		RECT	15.575 353.135 15.625 353.265 ;
		RECT	20.495 350.715 20.545 350.845 ;
		RECT	20.495 353.135 20.545 353.265 ;
		RECT	15.775 350.715 15.825 350.845 ;
		RECT	15.775 353.135 15.825 353.265 ;
		RECT	20.295 350.715 20.345 350.845 ;
		RECT	20.295 353.135 20.345 353.265 ;
		RECT	15.375 353.825 15.425 353.955 ;
		RECT	20.695 353.825 20.745 353.955 ;
		RECT	15.575 353.595 15.625 353.725 ;
		RECT	15.575 356.015 15.625 356.145 ;
		RECT	20.495 353.595 20.545 353.725 ;
		RECT	20.495 356.015 20.545 356.145 ;
		RECT	15.775 353.595 15.825 353.725 ;
		RECT	15.775 356.015 15.825 356.145 ;
		RECT	20.295 353.595 20.345 353.725 ;
		RECT	20.295 356.015 20.345 356.145 ;
		RECT	15.375 356.705 15.425 356.835 ;
		RECT	20.695 356.705 20.745 356.835 ;
		RECT	15.575 356.475 15.625 356.605 ;
		RECT	15.575 358.895 15.625 359.025 ;
		RECT	20.495 356.475 20.545 356.605 ;
		RECT	20.495 358.895 20.545 359.025 ;
		RECT	15.775 356.475 15.825 356.605 ;
		RECT	15.775 358.895 15.825 359.025 ;
		RECT	20.295 356.475 20.345 356.605 ;
		RECT	20.295 358.895 20.345 359.025 ;
		RECT	15.375 359.585 15.425 359.715 ;
		RECT	20.695 359.585 20.745 359.715 ;
		RECT	15.575 359.355 15.625 359.485 ;
		RECT	15.575 361.775 15.625 361.905 ;
		RECT	20.495 359.355 20.545 359.485 ;
		RECT	20.495 361.775 20.545 361.905 ;
		RECT	15.775 359.355 15.825 359.485 ;
		RECT	15.775 361.775 15.825 361.905 ;
		RECT	20.295 359.355 20.345 359.485 ;
		RECT	20.295 361.775 20.345 361.905 ;
		RECT	15.375 362.465 15.425 362.595 ;
		RECT	20.695 362.465 20.745 362.595 ;
		RECT	15.575 362.235 15.625 362.365 ;
		RECT	15.575 364.655 15.625 364.785 ;
		RECT	20.495 362.235 20.545 362.365 ;
		RECT	20.495 364.655 20.545 364.785 ;
		RECT	15.775 362.235 15.825 362.365 ;
		RECT	15.775 364.655 15.825 364.785 ;
		RECT	20.295 362.235 20.345 362.365 ;
		RECT	20.295 364.655 20.345 364.785 ;
		RECT	15.375 365.345 15.425 365.475 ;
		RECT	20.695 365.345 20.745 365.475 ;
		RECT	15.575 365.115 15.625 365.245 ;
		RECT	15.575 367.535 15.625 367.665 ;
		RECT	20.495 365.115 20.545 365.245 ;
		RECT	20.495 367.535 20.545 367.665 ;
		RECT	15.775 365.115 15.825 365.245 ;
		RECT	15.775 367.535 15.825 367.665 ;
		RECT	20.295 365.115 20.345 365.245 ;
		RECT	20.295 367.535 20.345 367.665 ;
		RECT	15.375 368.225 15.425 368.355 ;
		RECT	20.695 368.225 20.745 368.355 ;
		RECT	15.575 367.995 15.625 368.125 ;
		RECT	15.575 370.415 15.625 370.545 ;
		RECT	20.495 367.995 20.545 368.125 ;
		RECT	20.495 370.415 20.545 370.545 ;
		RECT	15.775 367.995 15.825 368.125 ;
		RECT	15.775 370.415 15.825 370.545 ;
		RECT	20.295 367.995 20.345 368.125 ;
		RECT	20.295 370.415 20.345 370.545 ;
		RECT	15.375 371.105 15.425 371.235 ;
		RECT	20.695 371.105 20.745 371.235 ;
		RECT	15.575 370.875 15.625 371.005 ;
		RECT	15.575 373.295 15.625 373.425 ;
		RECT	20.495 370.875 20.545 371.005 ;
		RECT	20.495 373.295 20.545 373.425 ;
		RECT	15.775 370.875 15.825 371.005 ;
		RECT	15.775 373.295 15.825 373.425 ;
		RECT	20.295 370.875 20.345 371.005 ;
		RECT	20.295 373.295 20.345 373.425 ;
		RECT	15.375 244.385 15.425 244.515 ;
		RECT	20.695 244.385 20.745 244.515 ;
		RECT	15.575 244.155 15.625 244.285 ;
		RECT	15.575 246.575 15.625 246.705 ;
		RECT	20.495 244.155 20.545 244.285 ;
		RECT	20.495 246.575 20.545 246.705 ;
		RECT	15.775 244.155 15.825 244.285 ;
		RECT	15.775 246.575 15.825 246.705 ;
		RECT	20.295 244.155 20.345 244.285 ;
		RECT	20.295 246.575 20.345 246.705 ;
		RECT	15.375 373.985 15.425 374.115 ;
		RECT	20.695 373.985 20.745 374.115 ;
		RECT	15.575 373.755 15.625 373.885 ;
		RECT	15.575 376.175 15.625 376.305 ;
		RECT	20.495 373.755 20.545 373.885 ;
		RECT	20.495 376.175 20.545 376.305 ;
		RECT	15.775 373.755 15.825 373.885 ;
		RECT	15.775 376.175 15.825 376.305 ;
		RECT	20.295 373.755 20.345 373.885 ;
		RECT	20.295 376.175 20.345 376.305 ;
		RECT	15.375 376.865 15.425 376.995 ;
		RECT	20.695 376.865 20.745 376.995 ;
		RECT	15.575 376.635 15.625 376.765 ;
		RECT	15.575 379.055 15.625 379.185 ;
		RECT	20.495 376.635 20.545 376.765 ;
		RECT	20.495 379.055 20.545 379.185 ;
		RECT	15.775 376.635 15.825 376.765 ;
		RECT	15.775 379.055 15.825 379.185 ;
		RECT	20.295 376.635 20.345 376.765 ;
		RECT	20.295 379.055 20.345 379.185 ;
		RECT	15.375 379.745 15.425 379.875 ;
		RECT	20.695 379.745 20.745 379.875 ;
		RECT	15.575 379.515 15.625 379.645 ;
		RECT	15.575 381.935 15.625 382.065 ;
		RECT	20.495 379.515 20.545 379.645 ;
		RECT	20.495 381.935 20.545 382.065 ;
		RECT	15.775 379.515 15.825 379.645 ;
		RECT	15.775 381.935 15.825 382.065 ;
		RECT	20.295 379.515 20.345 379.645 ;
		RECT	20.295 381.935 20.345 382.065 ;
		RECT	15.375 382.625 15.425 382.755 ;
		RECT	20.695 382.625 20.745 382.755 ;
		RECT	15.575 382.395 15.625 382.525 ;
		RECT	15.575 384.815 15.625 384.945 ;
		RECT	20.495 382.395 20.545 382.525 ;
		RECT	20.495 384.815 20.545 384.945 ;
		RECT	15.775 382.395 15.825 382.525 ;
		RECT	15.775 384.815 15.825 384.945 ;
		RECT	20.295 382.395 20.345 382.525 ;
		RECT	20.295 384.815 20.345 384.945 ;
		RECT	15.375 385.505 15.425 385.635 ;
		RECT	20.695 385.505 20.745 385.635 ;
		RECT	15.575 385.275 15.625 385.405 ;
		RECT	15.575 387.695 15.625 387.825 ;
		RECT	20.495 385.275 20.545 385.405 ;
		RECT	20.495 387.695 20.545 387.825 ;
		RECT	15.775 385.275 15.825 385.405 ;
		RECT	15.775 387.695 15.825 387.825 ;
		RECT	20.295 385.275 20.345 385.405 ;
		RECT	20.295 387.695 20.345 387.825 ;
		RECT	15.375 388.385 15.425 388.515 ;
		RECT	20.695 388.385 20.745 388.515 ;
		RECT	15.575 388.155 15.625 388.285 ;
		RECT	15.575 390.575 15.625 390.705 ;
		RECT	20.495 388.155 20.545 388.285 ;
		RECT	20.495 390.575 20.545 390.705 ;
		RECT	15.775 388.155 15.825 388.285 ;
		RECT	15.775 390.575 15.825 390.705 ;
		RECT	20.295 388.155 20.345 388.285 ;
		RECT	20.295 390.575 20.345 390.705 ;
		RECT	15.375 391.265 15.425 391.395 ;
		RECT	20.695 391.265 20.745 391.395 ;
		RECT	15.575 391.035 15.625 391.165 ;
		RECT	15.575 393.455 15.625 393.585 ;
		RECT	20.495 391.035 20.545 391.165 ;
		RECT	20.495 393.455 20.545 393.585 ;
		RECT	15.775 391.035 15.825 391.165 ;
		RECT	15.775 393.455 15.825 393.585 ;
		RECT	20.295 391.035 20.345 391.165 ;
		RECT	20.295 393.455 20.345 393.585 ;
		RECT	15.375 394.145 15.425 394.275 ;
		RECT	20.695 394.145 20.745 394.275 ;
		RECT	15.575 393.915 15.625 394.045 ;
		RECT	15.575 396.335 15.625 396.465 ;
		RECT	20.495 393.915 20.545 394.045 ;
		RECT	20.495 396.335 20.545 396.465 ;
		RECT	15.775 393.915 15.825 394.045 ;
		RECT	15.775 396.335 15.825 396.465 ;
		RECT	20.295 393.915 20.345 394.045 ;
		RECT	20.295 396.335 20.345 396.465 ;
		RECT	15.375 397.025 15.425 397.155 ;
		RECT	20.695 397.025 20.745 397.155 ;
		RECT	15.575 396.795 15.625 396.925 ;
		RECT	15.575 399.215 15.625 399.345 ;
		RECT	20.495 396.795 20.545 396.925 ;
		RECT	20.495 399.215 20.545 399.345 ;
		RECT	15.775 396.795 15.825 396.925 ;
		RECT	15.775 399.215 15.825 399.345 ;
		RECT	20.295 396.795 20.345 396.925 ;
		RECT	20.295 399.215 20.345 399.345 ;
		RECT	15.375 399.905 15.425 400.035 ;
		RECT	20.695 399.905 20.745 400.035 ;
		RECT	15.575 399.675 15.625 399.805 ;
		RECT	15.575 402.095 15.625 402.225 ;
		RECT	20.495 399.675 20.545 399.805 ;
		RECT	20.495 402.095 20.545 402.225 ;
		RECT	15.775 399.675 15.825 399.805 ;
		RECT	15.775 402.095 15.825 402.225 ;
		RECT	20.295 399.675 20.345 399.805 ;
		RECT	20.295 402.095 20.345 402.225 ;
		RECT	15.375 247.265 15.425 247.395 ;
		RECT	20.695 247.265 20.745 247.395 ;
		RECT	15.575 247.035 15.625 247.165 ;
		RECT	15.575 249.455 15.625 249.585 ;
		RECT	20.495 247.035 20.545 247.165 ;
		RECT	20.495 249.455 20.545 249.585 ;
		RECT	15.775 247.035 15.825 247.165 ;
		RECT	15.775 249.455 15.825 249.585 ;
		RECT	20.295 247.035 20.345 247.165 ;
		RECT	20.295 249.455 20.345 249.585 ;
		RECT	15.375 402.785 15.425 402.915 ;
		RECT	20.695 402.785 20.745 402.915 ;
		RECT	15.575 402.555 15.625 402.685 ;
		RECT	15.575 404.975 15.625 405.105 ;
		RECT	20.495 402.555 20.545 402.685 ;
		RECT	20.495 404.975 20.545 405.105 ;
		RECT	15.775 402.555 15.825 402.685 ;
		RECT	15.775 404.975 15.825 405.105 ;
		RECT	20.295 402.555 20.345 402.685 ;
		RECT	20.295 404.975 20.345 405.105 ;
		RECT	15.375 405.665 15.425 405.795 ;
		RECT	20.695 405.665 20.745 405.795 ;
		RECT	15.575 405.435 15.625 405.565 ;
		RECT	15.575 407.855 15.625 407.985 ;
		RECT	20.495 405.435 20.545 405.565 ;
		RECT	20.495 407.855 20.545 407.985 ;
		RECT	15.775 405.435 15.825 405.565 ;
		RECT	15.775 407.855 15.825 407.985 ;
		RECT	20.295 405.435 20.345 405.565 ;
		RECT	20.295 407.855 20.345 407.985 ;
		RECT	15.375 408.545 15.425 408.675 ;
		RECT	20.695 408.545 20.745 408.675 ;
		RECT	15.575 408.315 15.625 408.445 ;
		RECT	15.575 410.735 15.625 410.865 ;
		RECT	20.495 408.315 20.545 408.445 ;
		RECT	20.495 410.735 20.545 410.865 ;
		RECT	15.775 408.315 15.825 408.445 ;
		RECT	15.775 410.735 15.825 410.865 ;
		RECT	20.295 408.315 20.345 408.445 ;
		RECT	20.295 410.735 20.345 410.865 ;
		RECT	15.375 250.145 15.425 250.275 ;
		RECT	20.695 250.145 20.745 250.275 ;
		RECT	15.575 249.915 15.625 250.045 ;
		RECT	15.575 252.335 15.625 252.465 ;
		RECT	20.495 249.915 20.545 250.045 ;
		RECT	20.495 252.335 20.545 252.465 ;
		RECT	15.775 249.915 15.825 250.045 ;
		RECT	15.775 252.335 15.825 252.465 ;
		RECT	20.295 249.915 20.345 250.045 ;
		RECT	20.295 252.335 20.345 252.465 ;
		RECT	15.375 253.025 15.425 253.155 ;
		RECT	20.695 253.025 20.745 253.155 ;
		RECT	15.575 252.795 15.625 252.925 ;
		RECT	15.575 255.215 15.625 255.345 ;
		RECT	20.495 252.795 20.545 252.925 ;
		RECT	20.495 255.215 20.545 255.345 ;
		RECT	15.775 252.795 15.825 252.925 ;
		RECT	15.775 255.215 15.825 255.345 ;
		RECT	20.295 252.795 20.345 252.925 ;
		RECT	20.295 255.215 20.345 255.345 ;
		RECT	15.375 255.905 15.425 256.035 ;
		RECT	20.695 255.905 20.745 256.035 ;
		RECT	15.575 255.675 15.625 255.805 ;
		RECT	15.575 258.095 15.625 258.225 ;
		RECT	20.495 255.675 20.545 255.805 ;
		RECT	20.495 258.095 20.545 258.225 ;
		RECT	15.775 255.675 15.825 255.805 ;
		RECT	15.775 258.095 15.825 258.225 ;
		RECT	20.295 255.675 20.345 255.805 ;
		RECT	20.295 258.095 20.345 258.225 ;
		RECT	21.025 232.635 21.075 232.765 ;
		RECT	20.895 232.635 20.945 232.765 ;
		RECT	21.815 232.865 21.865 232.995 ;
		RECT	21.685 232.865 21.735 232.995 ;
		RECT	21.025 235.055 21.075 235.185 ;
		RECT	20.895 235.055 20.945 235.185 ;
		RECT	21.24 235.285 21.29 235.415 ;
		RECT	21.025 258.555 21.075 258.685 ;
		RECT	20.895 258.555 20.945 258.685 ;
		RECT	21.815 258.785 21.865 258.915 ;
		RECT	21.685 258.785 21.735 258.915 ;
		RECT	21.025 260.975 21.075 261.105 ;
		RECT	20.895 260.975 20.945 261.105 ;
		RECT	21.24 261.205 21.29 261.335 ;
		RECT	21.025 261.435 21.075 261.565 ;
		RECT	20.895 261.435 20.945 261.565 ;
		RECT	21.815 261.665 21.865 261.795 ;
		RECT	21.685 261.665 21.735 261.795 ;
		RECT	21.025 263.855 21.075 263.985 ;
		RECT	20.895 263.855 20.945 263.985 ;
		RECT	21.24 264.085 21.29 264.215 ;
		RECT	21.025 264.315 21.075 264.445 ;
		RECT	20.895 264.315 20.945 264.445 ;
		RECT	21.815 264.545 21.865 264.675 ;
		RECT	21.685 264.545 21.735 264.675 ;
		RECT	21.025 266.735 21.075 266.865 ;
		RECT	20.895 266.735 20.945 266.865 ;
		RECT	21.24 266.965 21.29 267.095 ;
		RECT	21.025 267.195 21.075 267.325 ;
		RECT	20.895 267.195 20.945 267.325 ;
		RECT	21.815 267.425 21.865 267.555 ;
		RECT	21.685 267.425 21.735 267.555 ;
		RECT	21.025 269.615 21.075 269.745 ;
		RECT	20.895 269.615 20.945 269.745 ;
		RECT	21.24 269.845 21.29 269.975 ;
		RECT	21.025 270.075 21.075 270.205 ;
		RECT	20.895 270.075 20.945 270.205 ;
		RECT	21.815 270.305 21.865 270.435 ;
		RECT	21.685 270.305 21.735 270.435 ;
		RECT	21.025 272.495 21.075 272.625 ;
		RECT	20.895 272.495 20.945 272.625 ;
		RECT	21.24 272.725 21.29 272.855 ;
		RECT	21.025 272.955 21.075 273.085 ;
		RECT	20.895 272.955 20.945 273.085 ;
		RECT	21.815 273.185 21.865 273.315 ;
		RECT	21.685 273.185 21.735 273.315 ;
		RECT	21.025 275.375 21.075 275.505 ;
		RECT	20.895 275.375 20.945 275.505 ;
		RECT	21.24 275.605 21.29 275.735 ;
		RECT	21.025 275.835 21.075 275.965 ;
		RECT	20.895 275.835 20.945 275.965 ;
		RECT	21.815 276.065 21.865 276.195 ;
		RECT	21.685 276.065 21.735 276.195 ;
		RECT	21.025 278.255 21.075 278.385 ;
		RECT	20.895 278.255 20.945 278.385 ;
		RECT	21.24 278.485 21.29 278.615 ;
		RECT	21.025 278.715 21.075 278.845 ;
		RECT	20.895 278.715 20.945 278.845 ;
		RECT	21.815 278.945 21.865 279.075 ;
		RECT	21.685 278.945 21.735 279.075 ;
		RECT	21.025 281.135 21.075 281.265 ;
		RECT	20.895 281.135 20.945 281.265 ;
		RECT	21.24 281.365 21.29 281.495 ;
		RECT	21.025 281.595 21.075 281.725 ;
		RECT	20.895 281.595 20.945 281.725 ;
		RECT	21.815 281.825 21.865 281.955 ;
		RECT	21.685 281.825 21.735 281.955 ;
		RECT	21.025 284.015 21.075 284.145 ;
		RECT	20.895 284.015 20.945 284.145 ;
		RECT	21.24 284.245 21.29 284.375 ;
		RECT	21.025 284.475 21.075 284.605 ;
		RECT	20.895 284.475 20.945 284.605 ;
		RECT	21.815 284.705 21.865 284.835 ;
		RECT	21.685 284.705 21.735 284.835 ;
		RECT	21.025 286.895 21.075 287.025 ;
		RECT	20.895 286.895 20.945 287.025 ;
		RECT	21.24 287.125 21.29 287.255 ;
		RECT	21.025 235.515 21.075 235.645 ;
		RECT	20.895 235.515 20.945 235.645 ;
		RECT	21.815 235.745 21.865 235.875 ;
		RECT	21.685 235.745 21.735 235.875 ;
		RECT	21.025 237.935 21.075 238.065 ;
		RECT	20.895 237.935 20.945 238.065 ;
		RECT	21.24 238.165 21.29 238.295 ;
		RECT	21.025 287.355 21.075 287.485 ;
		RECT	20.895 287.355 20.945 287.485 ;
		RECT	21.815 287.585 21.865 287.715 ;
		RECT	21.685 287.585 21.735 287.715 ;
		RECT	21.025 289.775 21.075 289.905 ;
		RECT	20.895 289.775 20.945 289.905 ;
		RECT	21.24 290.005 21.29 290.135 ;
		RECT	21.025 290.235 21.075 290.365 ;
		RECT	20.895 290.235 20.945 290.365 ;
		RECT	21.815 290.465 21.865 290.595 ;
		RECT	21.685 290.465 21.735 290.595 ;
		RECT	21.025 292.655 21.075 292.785 ;
		RECT	20.895 292.655 20.945 292.785 ;
		RECT	21.24 292.885 21.29 293.015 ;
		RECT	21.025 293.115 21.075 293.245 ;
		RECT	20.895 293.115 20.945 293.245 ;
		RECT	21.815 293.345 21.865 293.475 ;
		RECT	21.685 293.345 21.735 293.475 ;
		RECT	21.025 295.535 21.075 295.665 ;
		RECT	20.895 295.535 20.945 295.665 ;
		RECT	21.24 295.765 21.29 295.895 ;
		RECT	21.025 295.995 21.075 296.125 ;
		RECT	20.895 295.995 20.945 296.125 ;
		RECT	21.815 296.225 21.865 296.355 ;
		RECT	21.685 296.225 21.735 296.355 ;
		RECT	21.025 298.415 21.075 298.545 ;
		RECT	20.895 298.415 20.945 298.545 ;
		RECT	21.24 298.645 21.29 298.775 ;
		RECT	21.025 298.875 21.075 299.005 ;
		RECT	20.895 298.875 20.945 299.005 ;
		RECT	21.815 299.105 21.865 299.235 ;
		RECT	21.685 299.105 21.735 299.235 ;
		RECT	21.025 301.295 21.075 301.425 ;
		RECT	20.895 301.295 20.945 301.425 ;
		RECT	21.24 301.525 21.29 301.655 ;
		RECT	21.025 301.755 21.075 301.885 ;
		RECT	20.895 301.755 20.945 301.885 ;
		RECT	21.815 301.985 21.865 302.115 ;
		RECT	21.685 301.985 21.735 302.115 ;
		RECT	21.025 304.175 21.075 304.305 ;
		RECT	20.895 304.175 20.945 304.305 ;
		RECT	21.24 304.405 21.29 304.535 ;
		RECT	21.025 304.635 21.075 304.765 ;
		RECT	20.895 304.635 20.945 304.765 ;
		RECT	21.815 304.865 21.865 304.995 ;
		RECT	21.685 304.865 21.735 304.995 ;
		RECT	21.025 307.055 21.075 307.185 ;
		RECT	20.895 307.055 20.945 307.185 ;
		RECT	21.24 307.285 21.29 307.415 ;
		RECT	21.025 307.515 21.075 307.645 ;
		RECT	20.895 307.515 20.945 307.645 ;
		RECT	21.815 307.745 21.865 307.875 ;
		RECT	21.685 307.745 21.735 307.875 ;
		RECT	21.025 309.935 21.075 310.065 ;
		RECT	20.895 309.935 20.945 310.065 ;
		RECT	21.24 310.165 21.29 310.295 ;
		RECT	21.025 310.395 21.075 310.525 ;
		RECT	20.895 310.395 20.945 310.525 ;
		RECT	21.815 310.625 21.865 310.755 ;
		RECT	21.685 310.625 21.735 310.755 ;
		RECT	21.025 312.815 21.075 312.945 ;
		RECT	20.895 312.815 20.945 312.945 ;
		RECT	21.24 313.045 21.29 313.175 ;
		RECT	21.025 313.275 21.075 313.405 ;
		RECT	20.895 313.275 20.945 313.405 ;
		RECT	21.815 313.505 21.865 313.635 ;
		RECT	21.685 313.505 21.735 313.635 ;
		RECT	21.025 315.695 21.075 315.825 ;
		RECT	20.895 315.695 20.945 315.825 ;
		RECT	21.24 315.925 21.29 316.055 ;
		RECT	21.025 238.395 21.075 238.525 ;
		RECT	20.895 238.395 20.945 238.525 ;
		RECT	21.815 238.625 21.865 238.755 ;
		RECT	21.685 238.625 21.735 238.755 ;
		RECT	21.025 240.815 21.075 240.945 ;
		RECT	20.895 240.815 20.945 240.945 ;
		RECT	21.24 241.045 21.29 241.175 ;
		RECT	21.025 316.155 21.075 316.285 ;
		RECT	20.895 316.155 20.945 316.285 ;
		RECT	21.815 316.385 21.865 316.515 ;
		RECT	21.685 316.385 21.735 316.515 ;
		RECT	21.025 318.575 21.075 318.705 ;
		RECT	20.895 318.575 20.945 318.705 ;
		RECT	21.24 318.805 21.29 318.935 ;
		RECT	21.025 319.035 21.075 319.165 ;
		RECT	20.895 319.035 20.945 319.165 ;
		RECT	21.815 319.265 21.865 319.395 ;
		RECT	21.685 319.265 21.735 319.395 ;
		RECT	21.025 321.455 21.075 321.585 ;
		RECT	20.895 321.455 20.945 321.585 ;
		RECT	21.24 321.685 21.29 321.815 ;
		RECT	21.025 321.915 21.075 322.045 ;
		RECT	20.895 321.915 20.945 322.045 ;
		RECT	21.815 322.145 21.865 322.275 ;
		RECT	21.685 322.145 21.735 322.275 ;
		RECT	21.025 324.335 21.075 324.465 ;
		RECT	20.895 324.335 20.945 324.465 ;
		RECT	21.24 324.565 21.29 324.695 ;
		RECT	21.025 324.795 21.075 324.925 ;
		RECT	20.895 324.795 20.945 324.925 ;
		RECT	21.815 325.025 21.865 325.155 ;
		RECT	21.685 325.025 21.735 325.155 ;
		RECT	21.025 327.215 21.075 327.345 ;
		RECT	20.895 327.215 20.945 327.345 ;
		RECT	21.24 327.445 21.29 327.575 ;
		RECT	21.025 327.675 21.075 327.805 ;
		RECT	20.895 327.675 20.945 327.805 ;
		RECT	21.815 327.905 21.865 328.035 ;
		RECT	21.685 327.905 21.735 328.035 ;
		RECT	21.025 330.095 21.075 330.225 ;
		RECT	20.895 330.095 20.945 330.225 ;
		RECT	21.24 330.325 21.29 330.455 ;
		RECT	21.025 330.555 21.075 330.685 ;
		RECT	20.895 330.555 20.945 330.685 ;
		RECT	21.815 330.785 21.865 330.915 ;
		RECT	21.685 330.785 21.735 330.915 ;
		RECT	21.025 332.975 21.075 333.105 ;
		RECT	20.895 332.975 20.945 333.105 ;
		RECT	21.24 333.205 21.29 333.335 ;
		RECT	21.025 333.435 21.075 333.565 ;
		RECT	20.895 333.435 20.945 333.565 ;
		RECT	21.815 333.665 21.865 333.795 ;
		RECT	21.685 333.665 21.735 333.795 ;
		RECT	21.025 335.855 21.075 335.985 ;
		RECT	20.895 335.855 20.945 335.985 ;
		RECT	21.24 336.085 21.29 336.215 ;
		RECT	21.025 336.315 21.075 336.445 ;
		RECT	20.895 336.315 20.945 336.445 ;
		RECT	21.815 336.545 21.865 336.675 ;
		RECT	21.685 336.545 21.735 336.675 ;
		RECT	21.025 338.735 21.075 338.865 ;
		RECT	20.895 338.735 20.945 338.865 ;
		RECT	21.24 338.965 21.29 339.095 ;
		RECT	21.025 339.195 21.075 339.325 ;
		RECT	20.895 339.195 20.945 339.325 ;
		RECT	21.815 339.425 21.865 339.555 ;
		RECT	21.685 339.425 21.735 339.555 ;
		RECT	21.025 341.615 21.075 341.745 ;
		RECT	20.895 341.615 20.945 341.745 ;
		RECT	21.24 341.845 21.29 341.975 ;
		RECT	21.025 342.075 21.075 342.205 ;
		RECT	20.895 342.075 20.945 342.205 ;
		RECT	21.815 342.305 21.865 342.435 ;
		RECT	21.685 342.305 21.735 342.435 ;
		RECT	21.025 344.495 21.075 344.625 ;
		RECT	20.895 344.495 20.945 344.625 ;
		RECT	21.24 344.725 21.29 344.855 ;
		RECT	21.025 241.275 21.075 241.405 ;
		RECT	20.895 241.275 20.945 241.405 ;
		RECT	21.815 241.505 21.865 241.635 ;
		RECT	21.685 241.505 21.735 241.635 ;
		RECT	21.025 243.695 21.075 243.825 ;
		RECT	20.895 243.695 20.945 243.825 ;
		RECT	21.24 243.925 21.29 244.055 ;
		RECT	21.025 344.955 21.075 345.085 ;
		RECT	20.895 344.955 20.945 345.085 ;
		RECT	21.815 345.185 21.865 345.315 ;
		RECT	21.685 345.185 21.735 345.315 ;
		RECT	21.025 347.375 21.075 347.505 ;
		RECT	20.895 347.375 20.945 347.505 ;
		RECT	21.24 347.605 21.29 347.735 ;
		RECT	21.025 347.835 21.075 347.965 ;
		RECT	20.895 347.835 20.945 347.965 ;
		RECT	21.815 348.065 21.865 348.195 ;
		RECT	21.685 348.065 21.735 348.195 ;
		RECT	21.025 350.255 21.075 350.385 ;
		RECT	20.895 350.255 20.945 350.385 ;
		RECT	21.24 350.485 21.29 350.615 ;
		RECT	21.025 350.715 21.075 350.845 ;
		RECT	20.895 350.715 20.945 350.845 ;
		RECT	21.815 350.945 21.865 351.075 ;
		RECT	21.685 350.945 21.735 351.075 ;
		RECT	21.025 353.135 21.075 353.265 ;
		RECT	20.895 353.135 20.945 353.265 ;
		RECT	21.24 353.365 21.29 353.495 ;
		RECT	21.025 353.595 21.075 353.725 ;
		RECT	20.895 353.595 20.945 353.725 ;
		RECT	21.815 353.825 21.865 353.955 ;
		RECT	21.685 353.825 21.735 353.955 ;
		RECT	21.025 356.015 21.075 356.145 ;
		RECT	20.895 356.015 20.945 356.145 ;
		RECT	21.24 356.245 21.29 356.375 ;
		RECT	21.025 356.475 21.075 356.605 ;
		RECT	20.895 356.475 20.945 356.605 ;
		RECT	21.815 356.705 21.865 356.835 ;
		RECT	21.685 356.705 21.735 356.835 ;
		RECT	21.025 358.895 21.075 359.025 ;
		RECT	20.895 358.895 20.945 359.025 ;
		RECT	21.24 359.125 21.29 359.255 ;
		RECT	21.025 359.355 21.075 359.485 ;
		RECT	20.895 359.355 20.945 359.485 ;
		RECT	21.815 359.585 21.865 359.715 ;
		RECT	21.685 359.585 21.735 359.715 ;
		RECT	21.025 361.775 21.075 361.905 ;
		RECT	20.895 361.775 20.945 361.905 ;
		RECT	21.24 362.005 21.29 362.135 ;
		RECT	21.025 362.235 21.075 362.365 ;
		RECT	20.895 362.235 20.945 362.365 ;
		RECT	21.815 362.465 21.865 362.595 ;
		RECT	21.685 362.465 21.735 362.595 ;
		RECT	21.025 364.655 21.075 364.785 ;
		RECT	20.895 364.655 20.945 364.785 ;
		RECT	21.24 364.885 21.29 365.015 ;
		RECT	21.025 365.115 21.075 365.245 ;
		RECT	20.895 365.115 20.945 365.245 ;
		RECT	21.815 365.345 21.865 365.475 ;
		RECT	21.685 365.345 21.735 365.475 ;
		RECT	21.025 367.535 21.075 367.665 ;
		RECT	20.895 367.535 20.945 367.665 ;
		RECT	21.24 367.765 21.29 367.895 ;
		RECT	21.025 367.995 21.075 368.125 ;
		RECT	20.895 367.995 20.945 368.125 ;
		RECT	21.815 368.225 21.865 368.355 ;
		RECT	21.685 368.225 21.735 368.355 ;
		RECT	21.025 370.415 21.075 370.545 ;
		RECT	20.895 370.415 20.945 370.545 ;
		RECT	21.24 370.645 21.29 370.775 ;
		RECT	21.025 370.875 21.075 371.005 ;
		RECT	20.895 370.875 20.945 371.005 ;
		RECT	21.815 371.105 21.865 371.235 ;
		RECT	21.685 371.105 21.735 371.235 ;
		RECT	21.025 373.295 21.075 373.425 ;
		RECT	20.895 373.295 20.945 373.425 ;
		RECT	21.24 373.525 21.29 373.655 ;
		RECT	21.025 244.155 21.075 244.285 ;
		RECT	20.895 244.155 20.945 244.285 ;
		RECT	21.815 244.385 21.865 244.515 ;
		RECT	21.685 244.385 21.735 244.515 ;
		RECT	21.025 246.575 21.075 246.705 ;
		RECT	20.895 246.575 20.945 246.705 ;
		RECT	21.24 246.805 21.29 246.935 ;
		RECT	21.025 373.755 21.075 373.885 ;
		RECT	20.895 373.755 20.945 373.885 ;
		RECT	21.815 373.985 21.865 374.115 ;
		RECT	21.685 373.985 21.735 374.115 ;
		RECT	21.025 376.175 21.075 376.305 ;
		RECT	20.895 376.175 20.945 376.305 ;
		RECT	21.24 376.405 21.29 376.535 ;
		RECT	21.025 376.635 21.075 376.765 ;
		RECT	20.895 376.635 20.945 376.765 ;
		RECT	21.815 376.865 21.865 376.995 ;
		RECT	21.685 376.865 21.735 376.995 ;
		RECT	21.025 379.055 21.075 379.185 ;
		RECT	20.895 379.055 20.945 379.185 ;
		RECT	21.24 379.285 21.29 379.415 ;
		RECT	21.025 379.515 21.075 379.645 ;
		RECT	20.895 379.515 20.945 379.645 ;
		RECT	21.815 379.745 21.865 379.875 ;
		RECT	21.685 379.745 21.735 379.875 ;
		RECT	21.025 381.935 21.075 382.065 ;
		RECT	20.895 381.935 20.945 382.065 ;
		RECT	21.24 382.165 21.29 382.295 ;
		RECT	21.025 382.395 21.075 382.525 ;
		RECT	20.895 382.395 20.945 382.525 ;
		RECT	21.815 382.625 21.865 382.755 ;
		RECT	21.685 382.625 21.735 382.755 ;
		RECT	21.025 384.815 21.075 384.945 ;
		RECT	20.895 384.815 20.945 384.945 ;
		RECT	21.24 385.045 21.29 385.175 ;
		RECT	21.025 385.275 21.075 385.405 ;
		RECT	20.895 385.275 20.945 385.405 ;
		RECT	21.815 385.505 21.865 385.635 ;
		RECT	21.685 385.505 21.735 385.635 ;
		RECT	21.025 387.695 21.075 387.825 ;
		RECT	20.895 387.695 20.945 387.825 ;
		RECT	21.24 387.925 21.29 388.055 ;
		RECT	21.025 388.155 21.075 388.285 ;
		RECT	20.895 388.155 20.945 388.285 ;
		RECT	21.815 388.385 21.865 388.515 ;
		RECT	21.685 388.385 21.735 388.515 ;
		RECT	21.025 390.575 21.075 390.705 ;
		RECT	20.895 390.575 20.945 390.705 ;
		RECT	21.24 390.805 21.29 390.935 ;
		RECT	21.025 391.035 21.075 391.165 ;
		RECT	20.895 391.035 20.945 391.165 ;
		RECT	21.815 391.265 21.865 391.395 ;
		RECT	21.685 391.265 21.735 391.395 ;
		RECT	21.025 393.455 21.075 393.585 ;
		RECT	20.895 393.455 20.945 393.585 ;
		RECT	21.24 393.685 21.29 393.815 ;
		RECT	21.025 393.915 21.075 394.045 ;
		RECT	20.895 393.915 20.945 394.045 ;
		RECT	21.815 394.145 21.865 394.275 ;
		RECT	21.685 394.145 21.735 394.275 ;
		RECT	21.025 396.335 21.075 396.465 ;
		RECT	20.895 396.335 20.945 396.465 ;
		RECT	21.24 396.565 21.29 396.695 ;
		RECT	21.025 396.795 21.075 396.925 ;
		RECT	20.895 396.795 20.945 396.925 ;
		RECT	21.815 397.025 21.865 397.155 ;
		RECT	21.685 397.025 21.735 397.155 ;
		RECT	21.025 399.215 21.075 399.345 ;
		RECT	20.895 399.215 20.945 399.345 ;
		RECT	21.24 399.445 21.29 399.575 ;
		RECT	21.025 399.675 21.075 399.805 ;
		RECT	20.895 399.675 20.945 399.805 ;
		RECT	21.815 399.905 21.865 400.035 ;
		RECT	21.685 399.905 21.735 400.035 ;
		RECT	21.025 402.095 21.075 402.225 ;
		RECT	20.895 402.095 20.945 402.225 ;
		RECT	21.24 402.325 21.29 402.455 ;
		RECT	21.025 247.035 21.075 247.165 ;
		RECT	20.895 247.035 20.945 247.165 ;
		RECT	21.815 247.265 21.865 247.395 ;
		RECT	21.685 247.265 21.735 247.395 ;
		RECT	21.025 249.455 21.075 249.585 ;
		RECT	20.895 249.455 20.945 249.585 ;
		RECT	21.24 249.685 21.29 249.815 ;
		RECT	21.025 402.555 21.075 402.685 ;
		RECT	20.895 402.555 20.945 402.685 ;
		RECT	21.815 402.785 21.865 402.915 ;
		RECT	21.685 402.785 21.735 402.915 ;
		RECT	21.025 404.975 21.075 405.105 ;
		RECT	20.895 404.975 20.945 405.105 ;
		RECT	21.24 405.205 21.29 405.335 ;
		RECT	21.025 405.435 21.075 405.565 ;
		RECT	20.895 405.435 20.945 405.565 ;
		RECT	21.815 405.665 21.865 405.795 ;
		RECT	21.685 405.665 21.735 405.795 ;
		RECT	21.025 407.855 21.075 407.985 ;
		RECT	20.895 407.855 20.945 407.985 ;
		RECT	21.24 408.085 21.29 408.215 ;
		RECT	21.025 408.315 21.075 408.445 ;
		RECT	20.895 408.315 20.945 408.445 ;
		RECT	21.815 408.545 21.865 408.675 ;
		RECT	21.685 408.545 21.735 408.675 ;
		RECT	21.025 410.735 21.075 410.865 ;
		RECT	20.895 410.735 20.945 410.865 ;
		RECT	21.24 410.965 21.29 411.095 ;
		RECT	21.025 249.915 21.075 250.045 ;
		RECT	20.895 249.915 20.945 250.045 ;
		RECT	21.815 250.145 21.865 250.275 ;
		RECT	21.685 250.145 21.735 250.275 ;
		RECT	21.025 252.335 21.075 252.465 ;
		RECT	20.895 252.335 20.945 252.465 ;
		RECT	21.24 252.565 21.29 252.695 ;
		RECT	21.025 252.795 21.075 252.925 ;
		RECT	20.895 252.795 20.945 252.925 ;
		RECT	21.815 253.025 21.865 253.155 ;
		RECT	21.685 253.025 21.735 253.155 ;
		RECT	21.025 255.215 21.075 255.345 ;
		RECT	20.895 255.215 20.945 255.345 ;
		RECT	21.24 255.445 21.29 255.575 ;
		RECT	21.025 255.675 21.075 255.805 ;
		RECT	20.895 255.675 20.945 255.805 ;
		RECT	21.815 255.905 21.865 256.035 ;
		RECT	21.685 255.905 21.735 256.035 ;
		RECT	21.025 258.095 21.075 258.225 ;
		RECT	20.895 258.095 20.945 258.225 ;
		RECT	21.24 258.325 21.29 258.455 ;
		RECT	21.025 411.195 21.075 411.325 ;
		RECT	20.895 411.195 20.945 411.325 ;
		RECT	21.815 411.425 21.865 411.555 ;
		RECT	21.685 411.425 21.735 411.555 ;
		RECT	21.025 413.615 21.075 413.745 ;
		RECT	20.895 413.615 20.945 413.745 ;
		RECT	21.24 413.845 21.29 413.975 ;
		RECT	21.025 229.755 21.075 229.885 ;
		RECT	20.895 229.755 20.945 229.885 ;
		RECT	21.815 229.985 21.865 230.115 ;
		RECT	21.685 229.985 21.735 230.115 ;
		RECT	21.025 232.175 21.075 232.305 ;
		RECT	20.895 232.175 20.945 232.305 ;
		RECT	21.24 232.405 21.29 232.535 ;
		RECT	9.855 138.895 9.905 139.025 ;
		RECT	10.26 138.895 10.31 139.025 ;
		RECT	11.565 138.895 11.615 139.025 ;
		RECT	13.33 138.895 13.38 139.025 ;
		RECT	6.765 136.475 6.815 136.605 ;
		RECT	8.04 136.475 8.09 136.605 ;
		RECT	9.58 136.475 9.63 136.605 ;
		RECT	9.855 136.475 9.905 136.605 ;
		RECT	11.565 136.475 11.615 136.605 ;
		RECT	13.33 136.475 13.38 136.605 ;
		RECT	7.72 136.245 7.77 136.375 ;
		RECT	14.68 136.245 14.73 136.375 ;
		RECT	9.1 138.895 9.15 139.025 ;
		RECT	10.81 138.895 10.86 139.025 ;
		RECT	9.1 136.475 9.15 136.605 ;
		RECT	10.81 136.475 10.86 136.605 ;
		RECT	6.76 136.015 6.81 136.145 ;
		RECT	8.04 136.015 8.09 136.145 ;
		RECT	9.58 136.015 9.63 136.145 ;
		RECT	9.855 136.015 9.905 136.145 ;
		RECT	10.26 136.015 10.31 136.145 ;
		RECT	11.565 136.015 11.615 136.145 ;
		RECT	13.33 136.015 13.38 136.145 ;
		RECT	6.765 133.595 6.815 133.725 ;
		RECT	8.04 133.595 8.09 133.725 ;
		RECT	9.58 133.595 9.63 133.725 ;
		RECT	9.855 133.595 9.905 133.725 ;
		RECT	11.565 133.595 11.615 133.725 ;
		RECT	13.33 133.595 13.38 133.725 ;
		RECT	7.72 133.365 7.77 133.495 ;
		RECT	14.68 133.365 14.73 133.495 ;
		RECT	9.1 136.015 9.15 136.145 ;
		RECT	10.81 136.015 10.86 136.145 ;
		RECT	9.1 133.595 9.15 133.725 ;
		RECT	10.81 133.595 10.86 133.725 ;
		RECT	6.76 133.135 6.81 133.265 ;
		RECT	8.04 133.135 8.09 133.265 ;
		RECT	9.58 133.135 9.63 133.265 ;
		RECT	9.855 133.135 9.905 133.265 ;
		RECT	10.26 133.135 10.31 133.265 ;
		RECT	11.565 133.135 11.615 133.265 ;
		RECT	13.33 133.135 13.38 133.265 ;
		RECT	6.765 130.715 6.815 130.845 ;
		RECT	8.04 130.715 8.09 130.845 ;
		RECT	9.58 130.715 9.63 130.845 ;
		RECT	9.855 130.715 9.905 130.845 ;
		RECT	11.565 130.715 11.615 130.845 ;
		RECT	13.33 130.715 13.38 130.845 ;
		RECT	7.72 130.485 7.77 130.615 ;
		RECT	14.68 130.485 14.73 130.615 ;
		RECT	9.1 133.135 9.15 133.265 ;
		RECT	10.81 133.135 10.86 133.265 ;
		RECT	9.1 130.715 9.15 130.845 ;
		RECT	10.81 130.715 10.86 130.845 ;
		RECT	6.76 130.255 6.81 130.385 ;
		RECT	8.04 130.255 8.09 130.385 ;
		RECT	9.58 130.255 9.63 130.385 ;
		RECT	9.855 130.255 9.905 130.385 ;
		RECT	10.26 130.255 10.31 130.385 ;
		RECT	11.565 130.255 11.615 130.385 ;
		RECT	13.33 130.255 13.38 130.385 ;
		RECT	6.765 127.835 6.815 127.965 ;
		RECT	8.04 127.835 8.09 127.965 ;
		RECT	9.58 127.835 9.63 127.965 ;
		RECT	9.855 127.835 9.905 127.965 ;
		RECT	11.565 127.835 11.615 127.965 ;
		RECT	13.33 127.835 13.38 127.965 ;
		RECT	7.72 127.605 7.77 127.735 ;
		RECT	14.68 127.605 14.73 127.735 ;
		RECT	9.1 130.255 9.15 130.385 ;
		RECT	10.81 130.255 10.86 130.385 ;
		RECT	9.1 127.835 9.15 127.965 ;
		RECT	10.81 127.835 10.86 127.965 ;
		RECT	6.76 127.375 6.81 127.505 ;
		RECT	8.04 127.375 8.09 127.505 ;
		RECT	9.58 127.375 9.63 127.505 ;
		RECT	9.855 127.375 9.905 127.505 ;
		RECT	10.26 127.375 10.31 127.505 ;
		RECT	11.565 127.375 11.615 127.505 ;
		RECT	13.33 127.375 13.38 127.505 ;
		RECT	6.765 124.955 6.815 125.085 ;
		RECT	8.04 124.955 8.09 125.085 ;
		RECT	9.58 124.955 9.63 125.085 ;
		RECT	9.855 124.955 9.905 125.085 ;
		RECT	11.565 124.955 11.615 125.085 ;
		RECT	13.33 124.955 13.38 125.085 ;
		RECT	7.72 124.725 7.77 124.855 ;
		RECT	14.68 124.725 14.73 124.855 ;
		RECT	9.1 127.375 9.15 127.505 ;
		RECT	10.81 127.375 10.86 127.505 ;
		RECT	9.1 124.955 9.15 125.085 ;
		RECT	10.81 124.955 10.86 125.085 ;
		RECT	6.76 124.495 6.81 124.625 ;
		RECT	8.04 124.495 8.09 124.625 ;
		RECT	9.58 124.495 9.63 124.625 ;
		RECT	9.855 124.495 9.905 124.625 ;
		RECT	10.26 124.495 10.31 124.625 ;
		RECT	11.565 124.495 11.615 124.625 ;
		RECT	13.33 124.495 13.38 124.625 ;
		RECT	6.765 122.075 6.815 122.205 ;
		RECT	8.04 122.075 8.09 122.205 ;
		RECT	9.58 122.075 9.63 122.205 ;
		RECT	9.855 122.075 9.905 122.205 ;
		RECT	11.565 122.075 11.615 122.205 ;
		RECT	13.33 122.075 13.38 122.205 ;
		RECT	7.72 121.845 7.77 121.975 ;
		RECT	14.68 121.845 14.73 121.975 ;
		RECT	9.1 124.495 9.15 124.625 ;
		RECT	10.81 124.495 10.86 124.625 ;
		RECT	9.1 122.075 9.15 122.205 ;
		RECT	10.81 122.075 10.86 122.205 ;
		RECT	6.76 121.615 6.81 121.745 ;
		RECT	8.04 121.615 8.09 121.745 ;
		RECT	9.58 121.615 9.63 121.745 ;
		RECT	9.855 121.615 9.905 121.745 ;
		RECT	10.26 121.615 10.31 121.745 ;
		RECT	11.565 121.615 11.615 121.745 ;
		RECT	13.33 121.615 13.38 121.745 ;
		RECT	6.765 119.195 6.815 119.325 ;
		RECT	8.04 119.195 8.09 119.325 ;
		RECT	9.58 119.195 9.63 119.325 ;
		RECT	9.855 119.195 9.905 119.325 ;
		RECT	11.565 119.195 11.615 119.325 ;
		RECT	13.33 119.195 13.38 119.325 ;
		RECT	7.72 118.965 7.77 119.095 ;
		RECT	14.68 118.965 14.73 119.095 ;
		RECT	9.1 121.615 9.15 121.745 ;
		RECT	10.81 121.615 10.86 121.745 ;
		RECT	9.1 119.195 9.15 119.325 ;
		RECT	10.81 119.195 10.86 119.325 ;
		RECT	6.76 118.735 6.81 118.865 ;
		RECT	8.04 118.735 8.09 118.865 ;
		RECT	9.58 118.735 9.63 118.865 ;
		RECT	9.855 118.735 9.905 118.865 ;
		RECT	10.26 118.735 10.31 118.865 ;
		RECT	11.565 118.735 11.615 118.865 ;
		RECT	13.33 118.735 13.38 118.865 ;
		RECT	6.765 116.315 6.815 116.445 ;
		RECT	8.04 116.315 8.09 116.445 ;
		RECT	9.58 116.315 9.63 116.445 ;
		RECT	9.855 116.315 9.905 116.445 ;
		RECT	11.565 116.315 11.615 116.445 ;
		RECT	13.33 116.315 13.38 116.445 ;
		RECT	7.72 116.085 7.77 116.215 ;
		RECT	14.68 116.085 14.73 116.215 ;
		RECT	9.1 118.735 9.15 118.865 ;
		RECT	10.81 118.735 10.86 118.865 ;
		RECT	9.1 116.315 9.15 116.445 ;
		RECT	10.81 116.315 10.86 116.445 ;
		RECT	6.76 115.855 6.81 115.985 ;
		RECT	8.04 115.855 8.09 115.985 ;
		RECT	9.58 115.855 9.63 115.985 ;
		RECT	9.855 115.855 9.905 115.985 ;
		RECT	10.26 115.855 10.31 115.985 ;
		RECT	11.565 115.855 11.615 115.985 ;
		RECT	13.33 115.855 13.38 115.985 ;
		RECT	6.765 113.435 6.815 113.565 ;
		RECT	8.04 113.435 8.09 113.565 ;
		RECT	9.58 113.435 9.63 113.565 ;
		RECT	9.855 113.435 9.905 113.565 ;
		RECT	11.565 113.435 11.615 113.565 ;
		RECT	13.33 113.435 13.38 113.565 ;
		RECT	7.72 113.205 7.77 113.335 ;
		RECT	14.68 113.205 14.73 113.335 ;
		RECT	9.1 115.855 9.15 115.985 ;
		RECT	10.81 115.855 10.86 115.985 ;
		RECT	9.1 113.435 9.15 113.565 ;
		RECT	10.81 113.435 10.86 113.565 ;
		RECT	6.76 112.975 6.81 113.105 ;
		RECT	8.04 112.975 8.09 113.105 ;
		RECT	9.58 112.975 9.63 113.105 ;
		RECT	9.855 112.975 9.905 113.105 ;
		RECT	10.26 112.975 10.31 113.105 ;
		RECT	11.565 112.975 11.615 113.105 ;
		RECT	13.33 112.975 13.38 113.105 ;
		RECT	6.765 110.555 6.815 110.685 ;
		RECT	8.04 110.555 8.09 110.685 ;
		RECT	9.58 110.555 9.63 110.685 ;
		RECT	9.855 110.555 9.905 110.685 ;
		RECT	11.565 110.555 11.615 110.685 ;
		RECT	13.33 110.555 13.38 110.685 ;
		RECT	7.72 110.325 7.77 110.455 ;
		RECT	14.68 110.325 14.73 110.455 ;
		RECT	9.1 112.975 9.15 113.105 ;
		RECT	10.81 112.975 10.86 113.105 ;
		RECT	9.1 110.555 9.15 110.685 ;
		RECT	10.81 110.555 10.86 110.685 ;
		RECT	6.76 110.095 6.81 110.225 ;
		RECT	8.04 110.095 8.09 110.225 ;
		RECT	9.58 110.095 9.63 110.225 ;
		RECT	9.855 110.095 9.905 110.225 ;
		RECT	10.26 110.095 10.31 110.225 ;
		RECT	11.565 110.095 11.615 110.225 ;
		RECT	13.33 110.095 13.38 110.225 ;
		RECT	6.765 107.675 6.815 107.805 ;
		RECT	8.04 107.675 8.09 107.805 ;
		RECT	9.58 107.675 9.63 107.805 ;
		RECT	9.855 107.675 9.905 107.805 ;
		RECT	11.565 107.675 11.615 107.805 ;
		RECT	13.33 107.675 13.38 107.805 ;
		RECT	7.72 107.445 7.77 107.575 ;
		RECT	14.68 107.445 14.73 107.575 ;
		RECT	9.1 110.095 9.15 110.225 ;
		RECT	10.81 110.095 10.86 110.225 ;
		RECT	9.1 107.675 9.15 107.805 ;
		RECT	10.81 107.675 10.86 107.805 ;
		RECT	6.76 107.215 6.81 107.345 ;
		RECT	8.04 107.215 8.09 107.345 ;
		RECT	9.58 107.215 9.63 107.345 ;
		RECT	9.855 107.215 9.905 107.345 ;
		RECT	10.26 107.215 10.31 107.345 ;
		RECT	11.565 107.215 11.615 107.345 ;
		RECT	13.33 107.215 13.38 107.345 ;
		RECT	6.765 104.795 6.815 104.925 ;
		RECT	8.04 104.795 8.09 104.925 ;
		RECT	9.58 104.795 9.63 104.925 ;
		RECT	9.855 104.795 9.905 104.925 ;
		RECT	11.565 104.795 11.615 104.925 ;
		RECT	13.33 104.795 13.38 104.925 ;
		RECT	7.72 104.565 7.77 104.695 ;
		RECT	14.68 104.565 14.73 104.695 ;
		RECT	9.1 107.215 9.15 107.345 ;
		RECT	10.81 107.215 10.86 107.345 ;
		RECT	9.1 104.795 9.15 104.925 ;
		RECT	10.81 104.795 10.86 104.925 ;
		RECT	6.76 104.335 6.81 104.465 ;
		RECT	8.04 104.335 8.09 104.465 ;
		RECT	9.58 104.335 9.63 104.465 ;
		RECT	9.855 104.335 9.905 104.465 ;
		RECT	10.26 104.335 10.31 104.465 ;
		RECT	11.565 104.335 11.615 104.465 ;
		RECT	13.33 104.335 13.38 104.465 ;
		RECT	6.765 101.915 6.815 102.045 ;
		RECT	8.04 101.915 8.09 102.045 ;
		RECT	9.58 101.915 9.63 102.045 ;
		RECT	9.855 101.915 9.905 102.045 ;
		RECT	11.565 101.915 11.615 102.045 ;
		RECT	13.33 101.915 13.38 102.045 ;
		RECT	7.72 101.685 7.77 101.815 ;
		RECT	14.68 101.685 14.73 101.815 ;
		RECT	9.1 104.335 9.15 104.465 ;
		RECT	10.81 104.335 10.86 104.465 ;
		RECT	9.1 101.915 9.15 102.045 ;
		RECT	10.81 101.915 10.86 102.045 ;
		RECT	6.76 101.455 6.81 101.585 ;
		RECT	8.04 101.455 8.09 101.585 ;
		RECT	9.58 101.455 9.63 101.585 ;
		RECT	9.855 101.455 9.905 101.585 ;
		RECT	10.26 101.455 10.31 101.585 ;
		RECT	11.565 101.455 11.615 101.585 ;
		RECT	13.33 101.455 13.38 101.585 ;
		RECT	6.765 99.035 6.815 99.165 ;
		RECT	8.04 99.035 8.09 99.165 ;
		RECT	9.58 99.035 9.63 99.165 ;
		RECT	9.855 99.035 9.905 99.165 ;
		RECT	11.565 99.035 11.615 99.165 ;
		RECT	13.33 99.035 13.38 99.165 ;
		RECT	7.72 98.805 7.77 98.935 ;
		RECT	14.68 98.805 14.73 98.935 ;
		RECT	9.1 101.455 9.15 101.585 ;
		RECT	10.81 101.455 10.86 101.585 ;
		RECT	9.1 99.035 9.15 99.165 ;
		RECT	10.81 99.035 10.86 99.165 ;
		RECT	6.76 98.575 6.81 98.705 ;
		RECT	8.04 98.575 8.09 98.705 ;
		RECT	9.58 98.575 9.63 98.705 ;
		RECT	9.855 98.575 9.905 98.705 ;
		RECT	10.26 98.575 10.31 98.705 ;
		RECT	11.565 98.575 11.615 98.705 ;
		RECT	13.33 98.575 13.38 98.705 ;
		RECT	6.765 96.155 6.815 96.285 ;
		RECT	8.04 96.155 8.09 96.285 ;
		RECT	9.58 96.155 9.63 96.285 ;
		RECT	9.855 96.155 9.905 96.285 ;
		RECT	11.565 96.155 11.615 96.285 ;
		RECT	13.33 96.155 13.38 96.285 ;
		RECT	7.72 95.925 7.77 96.055 ;
		RECT	14.68 95.925 14.73 96.055 ;
		RECT	9.1 98.575 9.15 98.705 ;
		RECT	10.81 98.575 10.86 98.705 ;
		RECT	9.1 96.155 9.15 96.285 ;
		RECT	10.81 96.155 10.86 96.285 ;
		RECT	6.76 95.695 6.81 95.825 ;
		RECT	8.04 95.695 8.09 95.825 ;
		RECT	9.58 95.695 9.63 95.825 ;
		RECT	9.855 95.695 9.905 95.825 ;
		RECT	10.26 95.695 10.31 95.825 ;
		RECT	11.565 95.695 11.615 95.825 ;
		RECT	13.33 95.695 13.38 95.825 ;
		RECT	6.765 93.275 6.815 93.405 ;
		RECT	8.04 93.275 8.09 93.405 ;
		RECT	9.58 93.275 9.63 93.405 ;
		RECT	9.855 93.275 9.905 93.405 ;
		RECT	11.565 93.275 11.615 93.405 ;
		RECT	13.33 93.275 13.38 93.405 ;
		RECT	7.72 93.045 7.77 93.175 ;
		RECT	14.68 93.045 14.73 93.175 ;
		RECT	9.1 95.695 9.15 95.825 ;
		RECT	10.81 95.695 10.86 95.825 ;
		RECT	9.1 93.275 9.15 93.405 ;
		RECT	10.81 93.275 10.86 93.405 ;
		RECT	6.76 92.815 6.81 92.945 ;
		RECT	8.04 92.815 8.09 92.945 ;
		RECT	9.58 92.815 9.63 92.945 ;
		RECT	9.855 92.815 9.905 92.945 ;
		RECT	10.26 92.815 10.31 92.945 ;
		RECT	11.565 92.815 11.615 92.945 ;
		RECT	13.33 92.815 13.38 92.945 ;
		RECT	6.765 90.395 6.815 90.525 ;
		RECT	8.04 90.395 8.09 90.525 ;
		RECT	9.58 90.395 9.63 90.525 ;
		RECT	9.855 90.395 9.905 90.525 ;
		RECT	11.565 90.395 11.615 90.525 ;
		RECT	13.33 90.395 13.38 90.525 ;
		RECT	7.72 90.165 7.77 90.295 ;
		RECT	14.68 90.165 14.73 90.295 ;
		RECT	9.1 92.815 9.15 92.945 ;
		RECT	10.81 92.815 10.86 92.945 ;
		RECT	9.1 90.395 9.15 90.525 ;
		RECT	10.81 90.395 10.86 90.525 ;
		RECT	6.76 89.935 6.81 90.065 ;
		RECT	8.04 89.935 8.09 90.065 ;
		RECT	9.58 89.935 9.63 90.065 ;
		RECT	9.855 89.935 9.905 90.065 ;
		RECT	10.26 89.935 10.31 90.065 ;
		RECT	11.565 89.935 11.615 90.065 ;
		RECT	13.33 89.935 13.38 90.065 ;
		RECT	6.765 87.515 6.815 87.645 ;
		RECT	8.04 87.515 8.09 87.645 ;
		RECT	9.58 87.515 9.63 87.645 ;
		RECT	9.855 87.515 9.905 87.645 ;
		RECT	11.565 87.515 11.615 87.645 ;
		RECT	13.33 87.515 13.38 87.645 ;
		RECT	7.72 87.285 7.77 87.415 ;
		RECT	14.68 87.285 14.73 87.415 ;
		RECT	9.1 89.935 9.15 90.065 ;
		RECT	10.81 89.935 10.86 90.065 ;
		RECT	9.1 87.515 9.15 87.645 ;
		RECT	10.81 87.515 10.86 87.645 ;
		RECT	6.76 87.055 6.81 87.185 ;
		RECT	8.04 87.055 8.09 87.185 ;
		RECT	9.58 87.055 9.63 87.185 ;
		RECT	9.855 87.055 9.905 87.185 ;
		RECT	10.26 87.055 10.31 87.185 ;
		RECT	11.565 87.055 11.615 87.185 ;
		RECT	13.33 87.055 13.38 87.185 ;
		RECT	6.765 84.635 6.815 84.765 ;
		RECT	8.04 84.635 8.09 84.765 ;
		RECT	9.58 84.635 9.63 84.765 ;
		RECT	9.855 84.635 9.905 84.765 ;
		RECT	11.565 84.635 11.615 84.765 ;
		RECT	13.33 84.635 13.38 84.765 ;
		RECT	7.72 84.405 7.77 84.535 ;
		RECT	14.68 84.405 14.73 84.535 ;
		RECT	9.1 87.055 9.15 87.185 ;
		RECT	10.81 87.055 10.86 87.185 ;
		RECT	9.1 84.635 9.15 84.765 ;
		RECT	10.81 84.635 10.86 84.765 ;
		RECT	6.76 84.175 6.81 84.305 ;
		RECT	8.04 84.175 8.09 84.305 ;
		RECT	9.58 84.175 9.63 84.305 ;
		RECT	9.855 84.175 9.905 84.305 ;
		RECT	10.26 84.175 10.31 84.305 ;
		RECT	11.565 84.175 11.615 84.305 ;
		RECT	13.33 84.175 13.38 84.305 ;
		RECT	6.765 81.755 6.815 81.885 ;
		RECT	8.04 81.755 8.09 81.885 ;
		RECT	9.58 81.755 9.63 81.885 ;
		RECT	9.855 81.755 9.905 81.885 ;
		RECT	11.565 81.755 11.615 81.885 ;
		RECT	13.33 81.755 13.38 81.885 ;
		RECT	7.72 81.525 7.77 81.655 ;
		RECT	14.68 81.525 14.73 81.655 ;
		RECT	9.1 84.175 9.15 84.305 ;
		RECT	10.81 84.175 10.86 84.305 ;
		RECT	9.1 81.755 9.15 81.885 ;
		RECT	10.81 81.755 10.86 81.885 ;
		RECT	6.76 81.295 6.81 81.425 ;
		RECT	8.04 81.295 8.09 81.425 ;
		RECT	9.58 81.295 9.63 81.425 ;
		RECT	9.855 81.295 9.905 81.425 ;
		RECT	10.26 81.295 10.31 81.425 ;
		RECT	11.565 81.295 11.615 81.425 ;
		RECT	13.33 81.295 13.38 81.425 ;
		RECT	6.765 78.875 6.815 79.005 ;
		RECT	8.04 78.875 8.09 79.005 ;
		RECT	9.58 78.875 9.63 79.005 ;
		RECT	9.855 78.875 9.905 79.005 ;
		RECT	11.565 78.875 11.615 79.005 ;
		RECT	13.33 78.875 13.38 79.005 ;
		RECT	7.72 78.645 7.77 78.775 ;
		RECT	14.68 78.645 14.73 78.775 ;
		RECT	9.1 81.295 9.15 81.425 ;
		RECT	10.81 81.295 10.86 81.425 ;
		RECT	9.1 78.875 9.15 79.005 ;
		RECT	10.81 78.875 10.86 79.005 ;
		RECT	6.76 78.415 6.81 78.545 ;
		RECT	8.04 78.415 8.09 78.545 ;
		RECT	9.58 78.415 9.63 78.545 ;
		RECT	9.855 78.415 9.905 78.545 ;
		RECT	10.26 78.415 10.31 78.545 ;
		RECT	11.565 78.415 11.615 78.545 ;
		RECT	13.33 78.415 13.38 78.545 ;
		RECT	6.765 75.995 6.815 76.125 ;
		RECT	8.04 75.995 8.09 76.125 ;
		RECT	9.58 75.995 9.63 76.125 ;
		RECT	9.855 75.995 9.905 76.125 ;
		RECT	11.565 75.995 11.615 76.125 ;
		RECT	13.33 75.995 13.38 76.125 ;
		RECT	7.72 75.765 7.77 75.895 ;
		RECT	14.68 75.765 14.73 75.895 ;
		RECT	9.1 78.415 9.15 78.545 ;
		RECT	10.81 78.415 10.86 78.545 ;
		RECT	9.1 75.995 9.15 76.125 ;
		RECT	10.81 75.995 10.86 76.125 ;
		RECT	6.76 75.535 6.81 75.665 ;
		RECT	8.04 75.535 8.09 75.665 ;
		RECT	9.58 75.535 9.63 75.665 ;
		RECT	9.855 75.535 9.905 75.665 ;
		RECT	10.26 75.535 10.31 75.665 ;
		RECT	11.565 75.535 11.615 75.665 ;
		RECT	13.33 75.535 13.38 75.665 ;
		RECT	6.765 73.115 6.815 73.245 ;
		RECT	8.04 73.115 8.09 73.245 ;
		RECT	9.58 73.115 9.63 73.245 ;
		RECT	9.855 73.115 9.905 73.245 ;
		RECT	11.565 73.115 11.615 73.245 ;
		RECT	13.33 73.115 13.38 73.245 ;
		RECT	7.72 72.885 7.77 73.015 ;
		RECT	14.68 72.885 14.73 73.015 ;
		RECT	9.1 75.535 9.15 75.665 ;
		RECT	10.81 75.535 10.86 75.665 ;
		RECT	9.1 73.115 9.15 73.245 ;
		RECT	10.81 73.115 10.86 73.245 ;
		RECT	6.76 72.655 6.81 72.785 ;
		RECT	8.04 72.655 8.09 72.785 ;
		RECT	9.58 72.655 9.63 72.785 ;
		RECT	9.855 72.655 9.905 72.785 ;
		RECT	10.26 72.655 10.31 72.785 ;
		RECT	11.565 72.655 11.615 72.785 ;
		RECT	13.33 72.655 13.38 72.785 ;
		RECT	6.765 70.235 6.815 70.365 ;
		RECT	8.04 70.235 8.09 70.365 ;
		RECT	9.58 70.235 9.63 70.365 ;
		RECT	9.855 70.235 9.905 70.365 ;
		RECT	11.565 70.235 11.615 70.365 ;
		RECT	13.33 70.235 13.38 70.365 ;
		RECT	7.72 70.005 7.77 70.135 ;
		RECT	14.68 70.005 14.73 70.135 ;
		RECT	9.1 72.655 9.15 72.785 ;
		RECT	10.81 72.655 10.86 72.785 ;
		RECT	9.1 70.235 9.15 70.365 ;
		RECT	10.81 70.235 10.86 70.365 ;
		RECT	6.76 69.775 6.81 69.905 ;
		RECT	8.04 69.775 8.09 69.905 ;
		RECT	9.58 69.775 9.63 69.905 ;
		RECT	9.855 69.775 9.905 69.905 ;
		RECT	10.26 69.775 10.31 69.905 ;
		RECT	11.565 69.775 11.615 69.905 ;
		RECT	13.33 69.775 13.38 69.905 ;
		RECT	6.765 67.355 6.815 67.485 ;
		RECT	8.04 67.355 8.09 67.485 ;
		RECT	9.58 67.355 9.63 67.485 ;
		RECT	9.855 67.355 9.905 67.485 ;
		RECT	11.565 67.355 11.615 67.485 ;
		RECT	13.33 67.355 13.38 67.485 ;
		RECT	7.72 67.125 7.77 67.255 ;
		RECT	14.68 67.125 14.73 67.255 ;
		RECT	9.1 69.775 9.15 69.905 ;
		RECT	10.81 69.775 10.86 69.905 ;
		RECT	9.1 67.355 9.15 67.485 ;
		RECT	10.81 67.355 10.86 67.485 ;
		RECT	6.76 66.895 6.81 67.025 ;
		RECT	8.04 66.895 8.09 67.025 ;
		RECT	9.58 66.895 9.63 67.025 ;
		RECT	9.855 66.895 9.905 67.025 ;
		RECT	10.26 66.895 10.31 67.025 ;
		RECT	11.565 66.895 11.615 67.025 ;
		RECT	13.33 66.895 13.38 67.025 ;
		RECT	6.765 64.475 6.815 64.605 ;
		RECT	8.04 64.475 8.09 64.605 ;
		RECT	9.58 64.475 9.63 64.605 ;
		RECT	9.855 64.475 9.905 64.605 ;
		RECT	11.565 64.475 11.615 64.605 ;
		RECT	13.33 64.475 13.38 64.605 ;
		RECT	7.72 64.245 7.77 64.375 ;
		RECT	14.68 64.245 14.73 64.375 ;
		RECT	9.1 66.895 9.15 67.025 ;
		RECT	10.81 66.895 10.86 67.025 ;
		RECT	9.1 64.475 9.15 64.605 ;
		RECT	10.81 64.475 10.86 64.605 ;
		RECT	6.76 64.015 6.81 64.145 ;
		RECT	8.04 64.015 8.09 64.145 ;
		RECT	9.58 64.015 9.63 64.145 ;
		RECT	9.855 64.015 9.905 64.145 ;
		RECT	10.26 64.015 10.31 64.145 ;
		RECT	11.565 64.015 11.615 64.145 ;
		RECT	13.33 64.015 13.38 64.145 ;
		RECT	6.765 61.595 6.815 61.725 ;
		RECT	8.04 61.595 8.09 61.725 ;
		RECT	9.58 61.595 9.63 61.725 ;
		RECT	9.855 61.595 9.905 61.725 ;
		RECT	11.565 61.595 11.615 61.725 ;
		RECT	13.33 61.595 13.38 61.725 ;
		RECT	7.72 61.365 7.77 61.495 ;
		RECT	14.68 61.365 14.73 61.495 ;
		RECT	9.1 64.015 9.15 64.145 ;
		RECT	10.81 64.015 10.86 64.145 ;
		RECT	9.1 61.595 9.15 61.725 ;
		RECT	10.81 61.595 10.86 61.725 ;
		RECT	6.76 61.135 6.81 61.265 ;
		RECT	8.04 61.135 8.09 61.265 ;
		RECT	9.58 61.135 9.63 61.265 ;
		RECT	9.855 61.135 9.905 61.265 ;
		RECT	10.26 61.135 10.31 61.265 ;
		RECT	11.565 61.135 11.615 61.265 ;
		RECT	13.33 61.135 13.38 61.265 ;
		RECT	6.765 58.715 6.815 58.845 ;
		RECT	8.04 58.715 8.09 58.845 ;
		RECT	9.58 58.715 9.63 58.845 ;
		RECT	9.855 58.715 9.905 58.845 ;
		RECT	11.565 58.715 11.615 58.845 ;
		RECT	13.33 58.715 13.38 58.845 ;
		RECT	7.72 58.485 7.77 58.615 ;
		RECT	14.68 58.485 14.73 58.615 ;
		RECT	9.1 61.135 9.15 61.265 ;
		RECT	10.81 61.135 10.86 61.265 ;
		RECT	9.1 58.715 9.15 58.845 ;
		RECT	10.81 58.715 10.86 58.845 ;
		RECT	6.76 58.255 6.81 58.385 ;
		RECT	8.04 58.255 8.09 58.385 ;
		RECT	9.58 58.255 9.63 58.385 ;
		RECT	9.855 58.255 9.905 58.385 ;
		RECT	10.26 58.255 10.31 58.385 ;
		RECT	11.565 58.255 11.615 58.385 ;
		RECT	13.33 58.255 13.38 58.385 ;
		RECT	6.765 55.835 6.815 55.965 ;
		RECT	8.04 55.835 8.09 55.965 ;
		RECT	9.58 55.835 9.63 55.965 ;
		RECT	9.855 55.835 9.905 55.965 ;
		RECT	11.565 55.835 11.615 55.965 ;
		RECT	13.33 55.835 13.38 55.965 ;
		RECT	7.72 55.605 7.77 55.735 ;
		RECT	14.68 55.605 14.73 55.735 ;
		RECT	9.1 58.255 9.15 58.385 ;
		RECT	10.81 58.255 10.86 58.385 ;
		RECT	9.1 55.835 9.15 55.965 ;
		RECT	10.81 55.835 10.86 55.965 ;
		RECT	6.76 55.375 6.81 55.505 ;
		RECT	8.04 55.375 8.09 55.505 ;
		RECT	9.58 55.375 9.63 55.505 ;
		RECT	9.855 55.375 9.905 55.505 ;
		RECT	10.26 55.375 10.31 55.505 ;
		RECT	11.565 55.375 11.615 55.505 ;
		RECT	13.33 55.375 13.38 55.505 ;
		RECT	6.765 52.955 6.815 53.085 ;
		RECT	8.04 52.955 8.09 53.085 ;
		RECT	9.58 52.955 9.63 53.085 ;
		RECT	9.855 52.955 9.905 53.085 ;
		RECT	11.565 52.955 11.615 53.085 ;
		RECT	13.33 52.955 13.38 53.085 ;
		RECT	7.72 52.725 7.77 52.855 ;
		RECT	14.68 52.725 14.73 52.855 ;
		RECT	9.1 55.375 9.15 55.505 ;
		RECT	10.81 55.375 10.86 55.505 ;
		RECT	9.1 52.955 9.15 53.085 ;
		RECT	10.81 52.955 10.86 53.085 ;
		RECT	6.76 52.495 6.81 52.625 ;
		RECT	8.04 52.495 8.09 52.625 ;
		RECT	9.58 52.495 9.63 52.625 ;
		RECT	9.855 52.495 9.905 52.625 ;
		RECT	10.26 52.495 10.31 52.625 ;
		RECT	11.565 52.495 11.615 52.625 ;
		RECT	13.33 52.495 13.38 52.625 ;
		RECT	6.765 50.075 6.815 50.205 ;
		RECT	8.04 50.075 8.09 50.205 ;
		RECT	9.58 50.075 9.63 50.205 ;
		RECT	9.855 50.075 9.905 50.205 ;
		RECT	11.565 50.075 11.615 50.205 ;
		RECT	13.33 50.075 13.38 50.205 ;
		RECT	7.72 49.845 7.77 49.975 ;
		RECT	14.68 49.845 14.73 49.975 ;
		RECT	9.1 52.495 9.15 52.625 ;
		RECT	10.81 52.495 10.86 52.625 ;
		RECT	9.1 50.075 9.15 50.205 ;
		RECT	10.81 50.075 10.86 50.205 ;
		RECT	6.76 49.615 6.81 49.745 ;
		RECT	8.04 49.615 8.09 49.745 ;
		RECT	9.58 49.615 9.63 49.745 ;
		RECT	9.855 49.615 9.905 49.745 ;
		RECT	10.26 49.615 10.31 49.745 ;
		RECT	11.565 49.615 11.615 49.745 ;
		RECT	13.33 49.615 13.38 49.745 ;
		RECT	6.765 47.195 6.815 47.325 ;
		RECT	8.04 47.195 8.09 47.325 ;
		RECT	9.58 47.195 9.63 47.325 ;
		RECT	9.855 47.195 9.905 47.325 ;
		RECT	11.565 47.195 11.615 47.325 ;
		RECT	13.33 47.195 13.38 47.325 ;
		RECT	7.72 46.965 7.77 47.095 ;
		RECT	14.68 46.965 14.73 47.095 ;
		RECT	9.1 49.615 9.15 49.745 ;
		RECT	10.81 49.615 10.86 49.745 ;
		RECT	9.1 47.195 9.15 47.325 ;
		RECT	10.81 47.195 10.86 47.325 ;
		RECT	6.76 46.735 6.81 46.865 ;
		RECT	8.04 46.735 8.09 46.865 ;
		RECT	9.58 46.735 9.63 46.865 ;
		RECT	9.855 46.735 9.905 46.865 ;
		RECT	10.26 46.735 10.31 46.865 ;
		RECT	11.565 46.735 11.615 46.865 ;
		RECT	13.33 46.735 13.38 46.865 ;
		RECT	6.765 44.315 6.815 44.445 ;
		RECT	8.04 44.315 8.09 44.445 ;
		RECT	9.58 44.315 9.63 44.445 ;
		RECT	9.855 44.315 9.905 44.445 ;
		RECT	11.565 44.315 11.615 44.445 ;
		RECT	13.33 44.315 13.38 44.445 ;
		RECT	7.72 44.085 7.77 44.215 ;
		RECT	14.68 44.085 14.73 44.215 ;
		RECT	9.1 46.735 9.15 46.865 ;
		RECT	10.81 46.735 10.86 46.865 ;
		RECT	9.1 44.315 9.15 44.445 ;
		RECT	10.81 44.315 10.86 44.445 ;
		RECT	6.76 43.855 6.81 43.985 ;
		RECT	8.04 43.855 8.09 43.985 ;
		RECT	9.58 43.855 9.63 43.985 ;
		RECT	9.855 43.855 9.905 43.985 ;
		RECT	10.26 43.855 10.31 43.985 ;
		RECT	11.565 43.855 11.615 43.985 ;
		RECT	13.33 43.855 13.38 43.985 ;
		RECT	6.765 41.435 6.815 41.565 ;
		RECT	8.04 41.435 8.09 41.565 ;
		RECT	9.58 41.435 9.63 41.565 ;
		RECT	9.855 41.435 9.905 41.565 ;
		RECT	11.565 41.435 11.615 41.565 ;
		RECT	13.33 41.435 13.38 41.565 ;
		RECT	7.72 41.205 7.77 41.335 ;
		RECT	14.68 41.205 14.73 41.335 ;
		RECT	9.1 43.855 9.15 43.985 ;
		RECT	10.81 43.855 10.86 43.985 ;
		RECT	9.1 41.435 9.15 41.565 ;
		RECT	10.81 41.435 10.86 41.565 ;
		RECT	6.76 40.975 6.81 41.105 ;
		RECT	8.04 40.975 8.09 41.105 ;
		RECT	9.58 40.975 9.63 41.105 ;
		RECT	9.855 40.975 9.905 41.105 ;
		RECT	10.26 40.975 10.31 41.105 ;
		RECT	11.565 40.975 11.615 41.105 ;
		RECT	13.33 40.975 13.38 41.105 ;
		RECT	6.765 38.555 6.815 38.685 ;
		RECT	8.04 38.555 8.09 38.685 ;
		RECT	9.58 38.555 9.63 38.685 ;
		RECT	9.855 38.555 9.905 38.685 ;
		RECT	11.565 38.555 11.615 38.685 ;
		RECT	13.33 38.555 13.38 38.685 ;
		RECT	7.72 38.325 7.77 38.455 ;
		RECT	14.68 38.325 14.73 38.455 ;
		RECT	9.1 40.975 9.15 41.105 ;
		RECT	10.81 40.975 10.86 41.105 ;
		RECT	9.1 38.555 9.15 38.685 ;
		RECT	10.81 38.555 10.86 38.685 ;
		RECT	6.76 38.095 6.81 38.225 ;
		RECT	8.04 38.095 8.09 38.225 ;
		RECT	9.58 38.095 9.63 38.225 ;
		RECT	9.855 38.095 9.905 38.225 ;
		RECT	10.26 38.095 10.31 38.225 ;
		RECT	11.565 38.095 11.615 38.225 ;
		RECT	13.33 38.095 13.38 38.225 ;
		RECT	6.765 35.675 6.815 35.805 ;
		RECT	8.04 35.675 8.09 35.805 ;
		RECT	9.58 35.675 9.63 35.805 ;
		RECT	9.855 35.675 9.905 35.805 ;
		RECT	11.565 35.675 11.615 35.805 ;
		RECT	13.33 35.675 13.38 35.805 ;
		RECT	7.72 35.445 7.77 35.575 ;
		RECT	14.68 35.445 14.73 35.575 ;
		RECT	9.1 38.095 9.15 38.225 ;
		RECT	10.81 38.095 10.86 38.225 ;
		RECT	9.1 35.675 9.15 35.805 ;
		RECT	10.81 35.675 10.86 35.805 ;
		RECT	6.76 35.215 6.81 35.345 ;
		RECT	8.04 35.215 8.09 35.345 ;
		RECT	9.58 35.215 9.63 35.345 ;
		RECT	9.855 35.215 9.905 35.345 ;
		RECT	10.26 35.215 10.31 35.345 ;
		RECT	11.565 35.215 11.615 35.345 ;
		RECT	13.33 35.215 13.38 35.345 ;
		RECT	6.765 32.795 6.815 32.925 ;
		RECT	8.04 32.795 8.09 32.925 ;
		RECT	9.58 32.795 9.63 32.925 ;
		RECT	9.855 32.795 9.905 32.925 ;
		RECT	11.565 32.795 11.615 32.925 ;
		RECT	13.33 32.795 13.38 32.925 ;
		RECT	7.72 32.565 7.77 32.695 ;
		RECT	14.68 32.565 14.73 32.695 ;
		RECT	9.1 35.215 9.15 35.345 ;
		RECT	10.81 35.215 10.86 35.345 ;
		RECT	9.1 32.795 9.15 32.925 ;
		RECT	10.81 32.795 10.86 32.925 ;
		RECT	6.76 32.335 6.81 32.465 ;
		RECT	8.04 32.335 8.09 32.465 ;
		RECT	9.58 32.335 9.63 32.465 ;
		RECT	9.855 32.335 9.905 32.465 ;
		RECT	10.26 32.335 10.31 32.465 ;
		RECT	11.565 32.335 11.615 32.465 ;
		RECT	13.33 32.335 13.38 32.465 ;
		RECT	6.765 29.915 6.815 30.045 ;
		RECT	8.04 29.915 8.09 30.045 ;
		RECT	9.58 29.915 9.63 30.045 ;
		RECT	9.855 29.915 9.905 30.045 ;
		RECT	11.565 29.915 11.615 30.045 ;
		RECT	13.33 29.915 13.38 30.045 ;
		RECT	7.72 29.685 7.77 29.815 ;
		RECT	14.68 29.685 14.73 29.815 ;
		RECT	9.1 32.335 9.15 32.465 ;
		RECT	10.81 32.335 10.86 32.465 ;
		RECT	9.1 29.915 9.15 30.045 ;
		RECT	10.81 29.915 10.86 30.045 ;
		RECT	6.76 29.455 6.81 29.585 ;
		RECT	8.04 29.455 8.09 29.585 ;
		RECT	9.58 29.455 9.63 29.585 ;
		RECT	9.855 29.455 9.905 29.585 ;
		RECT	10.26 29.455 10.31 29.585 ;
		RECT	11.565 29.455 11.615 29.585 ;
		RECT	13.33 29.455 13.38 29.585 ;
		RECT	6.765 27.035 6.815 27.165 ;
		RECT	8.04 27.035 8.09 27.165 ;
		RECT	9.58 27.035 9.63 27.165 ;
		RECT	9.855 27.035 9.905 27.165 ;
		RECT	11.565 27.035 11.615 27.165 ;
		RECT	13.33 27.035 13.38 27.165 ;
		RECT	7.72 26.805 7.77 26.935 ;
		RECT	14.68 26.805 14.73 26.935 ;
		RECT	9.1 29.455 9.15 29.585 ;
		RECT	10.81 29.455 10.86 29.585 ;
		RECT	9.1 27.035 9.15 27.165 ;
		RECT	10.81 27.035 10.86 27.165 ;
		RECT	6.76 26.575 6.81 26.705 ;
		RECT	8.04 26.575 8.09 26.705 ;
		RECT	9.58 26.575 9.63 26.705 ;
		RECT	9.855 26.575 9.905 26.705 ;
		RECT	10.26 26.575 10.31 26.705 ;
		RECT	11.565 26.575 11.615 26.705 ;
		RECT	13.33 26.575 13.38 26.705 ;
		RECT	6.765 24.155 6.815 24.285 ;
		RECT	8.04 24.155 8.09 24.285 ;
		RECT	9.58 24.155 9.63 24.285 ;
		RECT	9.855 24.155 9.905 24.285 ;
		RECT	11.565 24.155 11.615 24.285 ;
		RECT	13.33 24.155 13.38 24.285 ;
		RECT	7.72 23.925 7.77 24.055 ;
		RECT	14.68 23.925 14.73 24.055 ;
		RECT	9.1 26.575 9.15 26.705 ;
		RECT	10.81 26.575 10.86 26.705 ;
		RECT	9.1 24.155 9.15 24.285 ;
		RECT	10.81 24.155 10.86 24.285 ;
		RECT	6.76 23.695 6.81 23.825 ;
		RECT	8.04 23.695 8.09 23.825 ;
		RECT	9.58 23.695 9.63 23.825 ;
		RECT	9.855 23.695 9.905 23.825 ;
		RECT	10.26 23.695 10.31 23.825 ;
		RECT	11.565 23.695 11.615 23.825 ;
		RECT	13.33 23.695 13.38 23.825 ;
		RECT	6.765 21.275 6.815 21.405 ;
		RECT	8.04 21.275 8.09 21.405 ;
		RECT	9.58 21.275 9.63 21.405 ;
		RECT	9.855 21.275 9.905 21.405 ;
		RECT	11.565 21.275 11.615 21.405 ;
		RECT	13.33 21.275 13.38 21.405 ;
		RECT	7.72 21.045 7.77 21.175 ;
		RECT	14.68 21.045 14.73 21.175 ;
		RECT	9.1 23.695 9.15 23.825 ;
		RECT	10.81 23.695 10.86 23.825 ;
		RECT	9.1 21.275 9.15 21.405 ;
		RECT	10.81 21.275 10.86 21.405 ;
		RECT	6.76 20.815 6.81 20.945 ;
		RECT	8.04 20.815 8.09 20.945 ;
		RECT	9.58 20.815 9.63 20.945 ;
		RECT	9.855 20.815 9.905 20.945 ;
		RECT	10.26 20.815 10.31 20.945 ;
		RECT	11.565 20.815 11.615 20.945 ;
		RECT	13.33 20.815 13.38 20.945 ;
		RECT	6.765 18.395 6.815 18.525 ;
		RECT	8.04 18.395 8.09 18.525 ;
		RECT	9.58 18.395 9.63 18.525 ;
		RECT	9.855 18.395 9.905 18.525 ;
		RECT	11.565 18.395 11.615 18.525 ;
		RECT	13.33 18.395 13.38 18.525 ;
		RECT	7.72 18.165 7.77 18.295 ;
		RECT	14.68 18.165 14.73 18.295 ;
		RECT	9.1 20.815 9.15 20.945 ;
		RECT	10.81 20.815 10.86 20.945 ;
		RECT	9.1 18.395 9.15 18.525 ;
		RECT	10.81 18.395 10.86 18.525 ;
		RECT	6.76 17.935 6.81 18.065 ;
		RECT	8.04 17.935 8.09 18.065 ;
		RECT	9.58 17.935 9.63 18.065 ;
		RECT	9.855 17.935 9.905 18.065 ;
		RECT	10.26 17.935 10.31 18.065 ;
		RECT	11.565 17.935 11.615 18.065 ;
		RECT	13.33 17.935 13.38 18.065 ;
		RECT	6.765 15.515 6.815 15.645 ;
		RECT	8.04 15.515 8.09 15.645 ;
		RECT	9.58 15.515 9.63 15.645 ;
		RECT	9.855 15.515 9.905 15.645 ;
		RECT	11.565 15.515 11.615 15.645 ;
		RECT	13.33 15.515 13.38 15.645 ;
		RECT	7.72 15.285 7.77 15.415 ;
		RECT	14.68 15.285 14.73 15.415 ;
		RECT	9.1 17.935 9.15 18.065 ;
		RECT	10.81 17.935 10.86 18.065 ;
		RECT	9.1 15.515 9.15 15.645 ;
		RECT	10.81 15.515 10.86 15.645 ;
		RECT	6.76 15.055 6.81 15.185 ;
		RECT	8.04 15.055 8.09 15.185 ;
		RECT	9.58 15.055 9.63 15.185 ;
		RECT	9.855 15.055 9.905 15.185 ;
		RECT	10.26 15.055 10.31 15.185 ;
		RECT	11.565 15.055 11.615 15.185 ;
		RECT	13.33 15.055 13.38 15.185 ;
		RECT	6.765 12.635 6.815 12.765 ;
		RECT	8.04 12.635 8.09 12.765 ;
		RECT	9.58 12.635 9.63 12.765 ;
		RECT	9.855 12.635 9.905 12.765 ;
		RECT	11.565 12.635 11.615 12.765 ;
		RECT	13.33 12.635 13.38 12.765 ;
		RECT	7.72 12.405 7.77 12.535 ;
		RECT	14.68 12.405 14.73 12.535 ;
		RECT	9.1 15.055 9.15 15.185 ;
		RECT	10.81 15.055 10.86 15.185 ;
		RECT	9.1 12.635 9.15 12.765 ;
		RECT	10.81 12.635 10.86 12.765 ;
		RECT	6.76 12.175 6.81 12.305 ;
		RECT	8.04 12.175 8.09 12.305 ;
		RECT	9.58 12.175 9.63 12.305 ;
		RECT	9.855 12.175 9.905 12.305 ;
		RECT	10.26 12.175 10.31 12.305 ;
		RECT	11.565 12.175 11.615 12.305 ;
		RECT	13.33 12.175 13.38 12.305 ;
		RECT	6.765 9.755 6.815 9.885 ;
		RECT	8.04 9.755 8.09 9.885 ;
		RECT	9.58 9.755 9.63 9.885 ;
		RECT	9.855 9.755 9.905 9.885 ;
		RECT	11.565 9.755 11.615 9.885 ;
		RECT	13.33 9.755 13.38 9.885 ;
		RECT	7.72 9.525 7.77 9.655 ;
		RECT	14.68 9.525 14.73 9.655 ;
		RECT	9.1 12.175 9.15 12.305 ;
		RECT	10.81 12.175 10.86 12.305 ;
		RECT	9.1 9.755 9.15 9.885 ;
		RECT	10.81 9.755 10.86 9.885 ;
		RECT	6.76 9.295 6.81 9.425 ;
		RECT	8.04 9.295 8.09 9.425 ;
		RECT	9.58 9.295 9.63 9.425 ;
		RECT	9.855 9.295 9.905 9.425 ;
		RECT	10.26 9.295 10.31 9.425 ;
		RECT	11.565 9.295 11.615 9.425 ;
		RECT	13.33 9.295 13.38 9.425 ;
		RECT	6.765 6.875 6.815 7.005 ;
		RECT	8.04 6.875 8.09 7.005 ;
		RECT	9.58 6.875 9.63 7.005 ;
		RECT	9.855 6.875 9.905 7.005 ;
		RECT	11.565 6.875 11.615 7.005 ;
		RECT	13.33 6.875 13.38 7.005 ;
		RECT	7.72 6.645 7.77 6.775 ;
		RECT	14.68 6.645 14.73 6.775 ;
		RECT	9.1 9.295 9.15 9.425 ;
		RECT	10.81 9.295 10.86 9.425 ;
		RECT	9.1 6.875 9.15 7.005 ;
		RECT	10.81 6.875 10.86 7.005 ;
		RECT	6.76 6.415 6.81 6.545 ;
		RECT	8.04 6.415 8.09 6.545 ;
		RECT	9.58 6.415 9.63 6.545 ;
		RECT	9.855 6.415 9.905 6.545 ;
		RECT	10.26 6.415 10.31 6.545 ;
		RECT	11.565 6.415 11.615 6.545 ;
		RECT	13.33 6.415 13.38 6.545 ;
		RECT	6.765 3.995 6.815 4.125 ;
		RECT	8.04 3.995 8.09 4.125 ;
		RECT	9.58 3.995 9.63 4.125 ;
		RECT	9.855 3.995 9.905 4.125 ;
		RECT	11.565 3.995 11.615 4.125 ;
		RECT	13.33 3.995 13.38 4.125 ;
		RECT	7.72 3.765 7.77 3.895 ;
		RECT	14.68 3.765 14.73 3.895 ;
		RECT	9.1 6.415 9.15 6.545 ;
		RECT	10.81 6.415 10.86 6.545 ;
		RECT	9.1 3.995 9.15 4.125 ;
		RECT	10.81 3.995 10.86 4.125 ;
		RECT	6.76 3.535 6.81 3.665 ;
		RECT	8.04 3.535 8.09 3.665 ;
		RECT	9.58 3.535 9.63 3.665 ;
		RECT	9.855 3.535 9.905 3.665 ;
		RECT	10.26 3.535 10.31 3.665 ;
		RECT	11.565 3.535 11.615 3.665 ;
		RECT	13.33 3.535 13.38 3.665 ;
		RECT	6.765 1.115 6.815 1.245 ;
		RECT	8.04 1.115 8.09 1.245 ;
		RECT	9.58 1.115 9.63 1.245 ;
		RECT	9.855 1.115 9.905 1.245 ;
		RECT	11.565 1.115 11.615 1.245 ;
		RECT	13.33 1.115 13.38 1.245 ;
		RECT	7.72 0.885 7.77 1.015 ;
		RECT	14.68 0.885 14.73 1.015 ;
		RECT	9.1 3.535 9.15 3.665 ;
		RECT	10.81 3.535 10.86 3.665 ;
		RECT	9.1 1.115 9.15 1.245 ;
		RECT	10.81 1.115 10.86 1.245 ;
		RECT	6.76 184.975 6.81 185.105 ;
		RECT	8.04 184.975 8.09 185.105 ;
		RECT	9.58 184.975 9.63 185.105 ;
		RECT	9.855 184.975 9.905 185.105 ;
		RECT	10.26 184.975 10.31 185.105 ;
		RECT	11.565 184.975 11.615 185.105 ;
		RECT	13.33 184.975 13.38 185.105 ;
		RECT	6.765 182.555 6.815 182.685 ;
		RECT	8.04 182.555 8.09 182.685 ;
		RECT	9.58 182.555 9.63 182.685 ;
		RECT	9.855 182.555 9.905 182.685 ;
		RECT	11.565 182.555 11.615 182.685 ;
		RECT	13.33 182.555 13.38 182.685 ;
		RECT	7.72 182.325 7.77 182.455 ;
		RECT	14.68 182.325 14.73 182.455 ;
		RECT	9.1 184.975 9.15 185.105 ;
		RECT	10.81 184.975 10.86 185.105 ;
		RECT	9.1 182.555 9.15 182.685 ;
		RECT	10.81 182.555 10.86 182.685 ;
		RECT	6.76 182.095 6.81 182.225 ;
		RECT	8.04 182.095 8.09 182.225 ;
		RECT	9.58 182.095 9.63 182.225 ;
		RECT	9.855 182.095 9.905 182.225 ;
		RECT	10.26 182.095 10.31 182.225 ;
		RECT	11.565 182.095 11.615 182.225 ;
		RECT	13.33 182.095 13.38 182.225 ;
		RECT	6.765 179.675 6.815 179.805 ;
		RECT	8.04 179.675 8.09 179.805 ;
		RECT	9.58 179.675 9.63 179.805 ;
		RECT	9.855 179.675 9.905 179.805 ;
		RECT	11.565 179.675 11.615 179.805 ;
		RECT	13.33 179.675 13.38 179.805 ;
		RECT	7.72 179.445 7.77 179.575 ;
		RECT	14.68 179.445 14.73 179.575 ;
		RECT	9.1 182.095 9.15 182.225 ;
		RECT	10.81 182.095 10.86 182.225 ;
		RECT	9.1 179.675 9.15 179.805 ;
		RECT	10.81 179.675 10.86 179.805 ;
		RECT	6.76 179.215 6.81 179.345 ;
		RECT	8.04 179.215 8.09 179.345 ;
		RECT	9.58 179.215 9.63 179.345 ;
		RECT	9.855 179.215 9.905 179.345 ;
		RECT	10.26 179.215 10.31 179.345 ;
		RECT	11.565 179.215 11.615 179.345 ;
		RECT	13.33 179.215 13.38 179.345 ;
		RECT	6.765 176.795 6.815 176.925 ;
		RECT	8.04 176.795 8.09 176.925 ;
		RECT	9.58 176.795 9.63 176.925 ;
		RECT	9.855 176.795 9.905 176.925 ;
		RECT	11.565 176.795 11.615 176.925 ;
		RECT	13.33 176.795 13.38 176.925 ;
		RECT	7.72 176.565 7.77 176.695 ;
		RECT	14.68 176.565 14.73 176.695 ;
		RECT	9.1 179.215 9.15 179.345 ;
		RECT	10.81 179.215 10.86 179.345 ;
		RECT	9.1 176.795 9.15 176.925 ;
		RECT	10.81 176.795 10.86 176.925 ;
		RECT	6.76 176.335 6.81 176.465 ;
		RECT	8.04 176.335 8.09 176.465 ;
		RECT	9.58 176.335 9.63 176.465 ;
		RECT	9.855 176.335 9.905 176.465 ;
		RECT	10.26 176.335 10.31 176.465 ;
		RECT	11.565 176.335 11.615 176.465 ;
		RECT	13.33 176.335 13.38 176.465 ;
		RECT	6.765 173.915 6.815 174.045 ;
		RECT	8.04 173.915 8.09 174.045 ;
		RECT	9.58 173.915 9.63 174.045 ;
		RECT	9.855 173.915 9.905 174.045 ;
		RECT	11.565 173.915 11.615 174.045 ;
		RECT	13.33 173.915 13.38 174.045 ;
		RECT	7.72 173.685 7.77 173.815 ;
		RECT	14.68 173.685 14.73 173.815 ;
		RECT	9.1 176.335 9.15 176.465 ;
		RECT	10.81 176.335 10.86 176.465 ;
		RECT	9.1 173.915 9.15 174.045 ;
		RECT	10.81 173.915 10.86 174.045 ;
		RECT	6.76 173.455 6.81 173.585 ;
		RECT	8.04 173.455 8.09 173.585 ;
		RECT	9.58 173.455 9.63 173.585 ;
		RECT	9.855 173.455 9.905 173.585 ;
		RECT	10.26 173.455 10.31 173.585 ;
		RECT	11.565 173.455 11.615 173.585 ;
		RECT	13.33 173.455 13.38 173.585 ;
		RECT	6.765 171.035 6.815 171.165 ;
		RECT	8.04 171.035 8.09 171.165 ;
		RECT	9.58 171.035 9.63 171.165 ;
		RECT	9.855 171.035 9.905 171.165 ;
		RECT	11.565 171.035 11.615 171.165 ;
		RECT	13.33 171.035 13.38 171.165 ;
		RECT	7.72 170.805 7.77 170.935 ;
		RECT	14.68 170.805 14.73 170.935 ;
		RECT	9.1 173.455 9.15 173.585 ;
		RECT	10.81 173.455 10.86 173.585 ;
		RECT	9.1 171.035 9.15 171.165 ;
		RECT	10.81 171.035 10.86 171.165 ;
		RECT	6.76 170.575 6.81 170.705 ;
		RECT	8.04 170.575 8.09 170.705 ;
		RECT	9.58 170.575 9.63 170.705 ;
		RECT	9.855 170.575 9.905 170.705 ;
		RECT	10.26 170.575 10.31 170.705 ;
		RECT	11.565 170.575 11.615 170.705 ;
		RECT	13.33 170.575 13.38 170.705 ;
		RECT	6.765 168.155 6.815 168.285 ;
		RECT	8.04 168.155 8.09 168.285 ;
		RECT	9.58 168.155 9.63 168.285 ;
		RECT	9.855 168.155 9.905 168.285 ;
		RECT	11.565 168.155 11.615 168.285 ;
		RECT	13.33 168.155 13.38 168.285 ;
		RECT	7.72 167.925 7.77 168.055 ;
		RECT	14.68 167.925 14.73 168.055 ;
		RECT	9.1 170.575 9.15 170.705 ;
		RECT	10.81 170.575 10.86 170.705 ;
		RECT	9.1 168.155 9.15 168.285 ;
		RECT	10.81 168.155 10.86 168.285 ;
		RECT	6.76 167.695 6.81 167.825 ;
		RECT	8.04 167.695 8.09 167.825 ;
		RECT	9.58 167.695 9.63 167.825 ;
		RECT	9.855 167.695 9.905 167.825 ;
		RECT	10.26 167.695 10.31 167.825 ;
		RECT	11.565 167.695 11.615 167.825 ;
		RECT	13.33 167.695 13.38 167.825 ;
		RECT	6.765 165.275 6.815 165.405 ;
		RECT	8.04 165.275 8.09 165.405 ;
		RECT	9.58 165.275 9.63 165.405 ;
		RECT	9.855 165.275 9.905 165.405 ;
		RECT	11.565 165.275 11.615 165.405 ;
		RECT	13.33 165.275 13.38 165.405 ;
		RECT	7.72 165.045 7.77 165.175 ;
		RECT	14.68 165.045 14.73 165.175 ;
		RECT	9.1 167.695 9.15 167.825 ;
		RECT	10.81 167.695 10.86 167.825 ;
		RECT	9.1 165.275 9.15 165.405 ;
		RECT	10.81 165.275 10.86 165.405 ;
		RECT	6.76 164.815 6.81 164.945 ;
		RECT	8.04 164.815 8.09 164.945 ;
		RECT	9.58 164.815 9.63 164.945 ;
		RECT	9.855 164.815 9.905 164.945 ;
		RECT	10.26 164.815 10.31 164.945 ;
		RECT	11.565 164.815 11.615 164.945 ;
		RECT	13.33 164.815 13.38 164.945 ;
		RECT	6.765 162.395 6.815 162.525 ;
		RECT	8.04 162.395 8.09 162.525 ;
		RECT	9.58 162.395 9.63 162.525 ;
		RECT	9.855 162.395 9.905 162.525 ;
		RECT	11.565 162.395 11.615 162.525 ;
		RECT	13.33 162.395 13.38 162.525 ;
		RECT	7.72 162.165 7.77 162.295 ;
		RECT	14.68 162.165 14.73 162.295 ;
		RECT	9.1 164.815 9.15 164.945 ;
		RECT	10.81 164.815 10.86 164.945 ;
		RECT	9.1 162.395 9.15 162.525 ;
		RECT	10.81 162.395 10.86 162.525 ;
		RECT	6.76 161.935 6.81 162.065 ;
		RECT	8.04 161.935 8.09 162.065 ;
		RECT	9.58 161.935 9.63 162.065 ;
		RECT	9.855 161.935 9.905 162.065 ;
		RECT	10.26 161.935 10.31 162.065 ;
		RECT	11.565 161.935 11.615 162.065 ;
		RECT	13.33 161.935 13.38 162.065 ;
		RECT	6.765 159.515 6.815 159.645 ;
		RECT	8.04 159.515 8.09 159.645 ;
		RECT	9.58 159.515 9.63 159.645 ;
		RECT	9.855 159.515 9.905 159.645 ;
		RECT	11.565 159.515 11.615 159.645 ;
		RECT	13.33 159.515 13.38 159.645 ;
		RECT	7.72 159.285 7.77 159.415 ;
		RECT	14.68 159.285 14.73 159.415 ;
		RECT	9.1 161.935 9.15 162.065 ;
		RECT	10.81 161.935 10.86 162.065 ;
		RECT	9.1 159.515 9.15 159.645 ;
		RECT	10.81 159.515 10.86 159.645 ;
		RECT	6.76 159.055 6.81 159.185 ;
		RECT	8.04 159.055 8.09 159.185 ;
		RECT	9.58 159.055 9.63 159.185 ;
		RECT	9.855 159.055 9.905 159.185 ;
		RECT	10.26 159.055 10.31 159.185 ;
		RECT	11.565 159.055 11.615 159.185 ;
		RECT	13.33 159.055 13.38 159.185 ;
		RECT	6.765 156.635 6.815 156.765 ;
		RECT	8.04 156.635 8.09 156.765 ;
		RECT	9.58 156.635 9.63 156.765 ;
		RECT	9.855 156.635 9.905 156.765 ;
		RECT	11.565 156.635 11.615 156.765 ;
		RECT	13.33 156.635 13.38 156.765 ;
		RECT	7.72 156.405 7.77 156.535 ;
		RECT	14.68 156.405 14.73 156.535 ;
		RECT	9.1 159.055 9.15 159.185 ;
		RECT	10.81 159.055 10.86 159.185 ;
		RECT	9.1 156.635 9.15 156.765 ;
		RECT	10.81 156.635 10.86 156.765 ;
		RECT	6.76 156.175 6.81 156.305 ;
		RECT	8.04 156.175 8.09 156.305 ;
		RECT	9.58 156.175 9.63 156.305 ;
		RECT	9.855 156.175 9.905 156.305 ;
		RECT	10.26 156.175 10.31 156.305 ;
		RECT	11.565 156.175 11.615 156.305 ;
		RECT	13.33 156.175 13.38 156.305 ;
		RECT	6.765 153.755 6.815 153.885 ;
		RECT	8.04 153.755 8.09 153.885 ;
		RECT	9.58 153.755 9.63 153.885 ;
		RECT	9.855 153.755 9.905 153.885 ;
		RECT	11.565 153.755 11.615 153.885 ;
		RECT	13.33 153.755 13.38 153.885 ;
		RECT	7.72 153.525 7.77 153.655 ;
		RECT	14.68 153.525 14.73 153.655 ;
		RECT	9.1 156.175 9.15 156.305 ;
		RECT	10.81 156.175 10.86 156.305 ;
		RECT	9.1 153.755 9.15 153.885 ;
		RECT	10.81 153.755 10.86 153.885 ;
		RECT	6.76 153.295 6.81 153.425 ;
		RECT	8.04 153.295 8.09 153.425 ;
		RECT	9.58 153.295 9.63 153.425 ;
		RECT	9.855 153.295 9.905 153.425 ;
		RECT	10.26 153.295 10.31 153.425 ;
		RECT	11.565 153.295 11.615 153.425 ;
		RECT	13.33 153.295 13.38 153.425 ;
		RECT	6.765 150.875 6.815 151.005 ;
		RECT	8.04 150.875 8.09 151.005 ;
		RECT	9.58 150.875 9.63 151.005 ;
		RECT	9.855 150.875 9.905 151.005 ;
		RECT	11.565 150.875 11.615 151.005 ;
		RECT	13.33 150.875 13.38 151.005 ;
		RECT	7.72 150.645 7.77 150.775 ;
		RECT	14.68 150.645 14.73 150.775 ;
		RECT	9.1 153.295 9.15 153.425 ;
		RECT	10.81 153.295 10.86 153.425 ;
		RECT	9.1 150.875 9.15 151.005 ;
		RECT	10.81 150.875 10.86 151.005 ;
		RECT	6.76 150.415 6.81 150.545 ;
		RECT	8.04 150.415 8.09 150.545 ;
		RECT	9.58 150.415 9.63 150.545 ;
		RECT	9.855 150.415 9.905 150.545 ;
		RECT	10.26 150.415 10.31 150.545 ;
		RECT	11.565 150.415 11.615 150.545 ;
		RECT	13.33 150.415 13.38 150.545 ;
		RECT	6.765 147.995 6.815 148.125 ;
		RECT	8.04 147.995 8.09 148.125 ;
		RECT	9.58 147.995 9.63 148.125 ;
		RECT	9.855 147.995 9.905 148.125 ;
		RECT	11.565 147.995 11.615 148.125 ;
		RECT	13.33 147.995 13.38 148.125 ;
		RECT	7.72 147.765 7.77 147.895 ;
		RECT	14.68 147.765 14.73 147.895 ;
		RECT	9.1 150.415 9.15 150.545 ;
		RECT	10.81 150.415 10.86 150.545 ;
		RECT	9.1 147.995 9.15 148.125 ;
		RECT	10.81 147.995 10.86 148.125 ;
		RECT	6.76 147.535 6.81 147.665 ;
		RECT	8.04 147.535 8.09 147.665 ;
		RECT	9.58 147.535 9.63 147.665 ;
		RECT	9.855 147.535 9.905 147.665 ;
		RECT	10.26 147.535 10.31 147.665 ;
		RECT	11.565 147.535 11.615 147.665 ;
		RECT	13.33 147.535 13.38 147.665 ;
		RECT	6.765 145.115 6.815 145.245 ;
		RECT	8.04 145.115 8.09 145.245 ;
		RECT	9.58 145.115 9.63 145.245 ;
		RECT	9.855 145.115 9.905 145.245 ;
		RECT	11.565 145.115 11.615 145.245 ;
		RECT	13.33 145.115 13.38 145.245 ;
		RECT	7.72 144.885 7.77 145.015 ;
		RECT	14.68 144.885 14.73 145.015 ;
		RECT	9.1 147.535 9.15 147.665 ;
		RECT	10.81 147.535 10.86 147.665 ;
		RECT	9.1 145.115 9.15 145.245 ;
		RECT	10.81 145.115 10.86 145.245 ;
		RECT	6.76 144.655 6.81 144.785 ;
		RECT	8.04 144.655 8.09 144.785 ;
		RECT	9.58 144.655 9.63 144.785 ;
		RECT	9.855 144.655 9.905 144.785 ;
		RECT	10.26 144.655 10.31 144.785 ;
		RECT	11.565 144.655 11.615 144.785 ;
		RECT	13.33 144.655 13.38 144.785 ;
		RECT	6.765 142.235 6.815 142.365 ;
		RECT	8.04 142.235 8.09 142.365 ;
		RECT	9.58 142.235 9.63 142.365 ;
		RECT	9.855 142.235 9.905 142.365 ;
		RECT	11.565 142.235 11.615 142.365 ;
		RECT	13.33 142.235 13.38 142.365 ;
		RECT	7.72 142.005 7.77 142.135 ;
		RECT	14.68 142.005 14.73 142.135 ;
		RECT	9.1 144.655 9.15 144.785 ;
		RECT	10.81 144.655 10.86 144.785 ;
		RECT	9.1 142.235 9.15 142.365 ;
		RECT	10.81 142.235 10.86 142.365 ;
		RECT	6.76 141.775 6.81 141.905 ;
		RECT	8.04 141.775 8.09 141.905 ;
		RECT	9.58 141.775 9.63 141.905 ;
		RECT	9.855 141.775 9.905 141.905 ;
		RECT	10.26 141.775 10.31 141.905 ;
		RECT	11.565 141.775 11.615 141.905 ;
		RECT	13.33 141.775 13.38 141.905 ;
		RECT	6.765 139.355 6.815 139.485 ;
		RECT	8.04 139.355 8.09 139.485 ;
		RECT	9.58 139.355 9.63 139.485 ;
		RECT	9.855 139.355 9.905 139.485 ;
		RECT	11.565 139.355 11.615 139.485 ;
		RECT	13.33 139.355 13.38 139.485 ;
		RECT	7.72 139.125 7.77 139.255 ;
		RECT	14.68 139.125 14.73 139.255 ;
		RECT	9.1 141.775 9.15 141.905 ;
		RECT	10.81 141.775 10.86 141.905 ;
		RECT	9.1 139.355 9.15 139.485 ;
		RECT	10.81 139.355 10.86 139.485 ;
		RECT	6.76 138.895 6.81 139.025 ;
		RECT	8.04 138.895 8.09 139.025 ;
		RECT	9.58 138.895 9.63 139.025 ;
		RECT	14.87 182.095 14.92 182.225 ;
		RECT	6.76 181.635 6.81 181.765 ;
		RECT	8.04 181.635 8.09 181.765 ;
		RECT	9.58 181.635 9.63 181.765 ;
		RECT	9.855 181.635 9.905 181.765 ;
		RECT	10.26 181.635 10.31 181.765 ;
		RECT	11.565 181.635 11.615 181.765 ;
		RECT	13.33 181.635 13.38 181.765 ;
		RECT	14.23 181.635 14.28 181.765 ;
		RECT	14.23 179.905 14.28 180.035 ;
		RECT	14.87 179.675 14.92 179.805 ;
		RECT	6.215 179.445 6.265 179.575 ;
		RECT	6.605 179.445 6.655 179.575 ;
		RECT	7.265 179.445 7.315 179.575 ;
		RECT	8.96 179.445 9.01 179.575 ;
		RECT	9.31 179.445 9.36 179.575 ;
		RECT	12.095 179.445 12.145 179.575 ;
		RECT	12.355 179.445 12.405 179.575 ;
		RECT	13.06 179.445 13.11 179.575 ;
		RECT	14.52 179.445 14.57 179.575 ;
		RECT	14.87 156.175 14.92 156.305 ;
		RECT	6.76 155.715 6.81 155.845 ;
		RECT	8.04 155.715 8.09 155.845 ;
		RECT	9.58 155.715 9.63 155.845 ;
		RECT	9.855 155.715 9.905 155.845 ;
		RECT	10.26 155.715 10.31 155.845 ;
		RECT	11.565 155.715 11.615 155.845 ;
		RECT	13.33 155.715 13.38 155.845 ;
		RECT	14.23 155.715 14.28 155.845 ;
		RECT	14.23 153.985 14.28 154.115 ;
		RECT	14.87 153.755 14.92 153.885 ;
		RECT	6.215 153.525 6.265 153.655 ;
		RECT	6.605 153.525 6.655 153.655 ;
		RECT	7.265 153.525 7.315 153.655 ;
		RECT	8.96 153.525 9.01 153.655 ;
		RECT	9.31 153.525 9.36 153.655 ;
		RECT	12.095 153.525 12.145 153.655 ;
		RECT	12.355 153.525 12.405 153.655 ;
		RECT	13.06 153.525 13.11 153.655 ;
		RECT	14.52 153.525 14.57 153.655 ;
		RECT	14.87 153.295 14.92 153.425 ;
		RECT	6.76 152.835 6.81 152.965 ;
		RECT	8.04 152.835 8.09 152.965 ;
		RECT	9.58 152.835 9.63 152.965 ;
		RECT	9.855 152.835 9.905 152.965 ;
		RECT	10.26 152.835 10.31 152.965 ;
		RECT	11.565 152.835 11.615 152.965 ;
		RECT	13.33 152.835 13.38 152.965 ;
		RECT	14.23 152.835 14.28 152.965 ;
		RECT	14.23 151.105 14.28 151.235 ;
		RECT	14.87 150.875 14.92 151.005 ;
		RECT	6.215 150.645 6.265 150.775 ;
		RECT	6.605 150.645 6.655 150.775 ;
		RECT	7.265 150.645 7.315 150.775 ;
		RECT	8.96 150.645 9.01 150.775 ;
		RECT	9.31 150.645 9.36 150.775 ;
		RECT	12.095 150.645 12.145 150.775 ;
		RECT	12.355 150.645 12.405 150.775 ;
		RECT	13.06 150.645 13.11 150.775 ;
		RECT	14.52 150.645 14.57 150.775 ;
		RECT	14.87 150.415 14.92 150.545 ;
		RECT	6.76 149.955 6.81 150.085 ;
		RECT	8.04 149.955 8.09 150.085 ;
		RECT	9.58 149.955 9.63 150.085 ;
		RECT	9.855 149.955 9.905 150.085 ;
		RECT	10.26 149.955 10.31 150.085 ;
		RECT	11.565 149.955 11.615 150.085 ;
		RECT	13.33 149.955 13.38 150.085 ;
		RECT	14.23 149.955 14.28 150.085 ;
		RECT	14.23 148.225 14.28 148.355 ;
		RECT	14.87 147.995 14.92 148.125 ;
		RECT	6.215 147.765 6.265 147.895 ;
		RECT	6.605 147.765 6.655 147.895 ;
		RECT	7.265 147.765 7.315 147.895 ;
		RECT	8.96 147.765 9.01 147.895 ;
		RECT	9.31 147.765 9.36 147.895 ;
		RECT	12.095 147.765 12.145 147.895 ;
		RECT	12.355 147.765 12.405 147.895 ;
		RECT	13.06 147.765 13.11 147.895 ;
		RECT	14.52 147.765 14.57 147.895 ;
		RECT	14.87 147.535 14.92 147.665 ;
		RECT	6.76 147.075 6.81 147.205 ;
		RECT	8.04 147.075 8.09 147.205 ;
		RECT	9.58 147.075 9.63 147.205 ;
		RECT	9.855 147.075 9.905 147.205 ;
		RECT	10.26 147.075 10.31 147.205 ;
		RECT	11.565 147.075 11.615 147.205 ;
		RECT	13.33 147.075 13.38 147.205 ;
		RECT	14.23 147.075 14.28 147.205 ;
		RECT	14.23 145.345 14.28 145.475 ;
		RECT	14.87 145.115 14.92 145.245 ;
		RECT	6.215 144.885 6.265 145.015 ;
		RECT	6.605 144.885 6.655 145.015 ;
		RECT	7.265 144.885 7.315 145.015 ;
		RECT	8.96 144.885 9.01 145.015 ;
		RECT	9.31 144.885 9.36 145.015 ;
		RECT	12.095 144.885 12.145 145.015 ;
		RECT	12.355 144.885 12.405 145.015 ;
		RECT	13.06 144.885 13.11 145.015 ;
		RECT	14.52 144.885 14.57 145.015 ;
		RECT	14.87 144.655 14.92 144.785 ;
		RECT	6.76 144.195 6.81 144.325 ;
		RECT	8.04 144.195 8.09 144.325 ;
		RECT	9.58 144.195 9.63 144.325 ;
		RECT	9.855 144.195 9.905 144.325 ;
		RECT	10.26 144.195 10.31 144.325 ;
		RECT	11.565 144.195 11.615 144.325 ;
		RECT	13.33 144.195 13.38 144.325 ;
		RECT	14.23 144.195 14.28 144.325 ;
		RECT	14.23 142.465 14.28 142.595 ;
		RECT	14.87 142.235 14.92 142.365 ;
		RECT	6.215 142.005 6.265 142.135 ;
		RECT	6.605 142.005 6.655 142.135 ;
		RECT	7.265 142.005 7.315 142.135 ;
		RECT	8.96 142.005 9.01 142.135 ;
		RECT	9.31 142.005 9.36 142.135 ;
		RECT	12.095 142.005 12.145 142.135 ;
		RECT	12.355 142.005 12.405 142.135 ;
		RECT	13.06 142.005 13.11 142.135 ;
		RECT	14.52 142.005 14.57 142.135 ;
		RECT	14.87 141.775 14.92 141.905 ;
		RECT	6.76 141.315 6.81 141.445 ;
		RECT	8.04 141.315 8.09 141.445 ;
		RECT	9.58 141.315 9.63 141.445 ;
		RECT	9.855 141.315 9.905 141.445 ;
		RECT	10.26 141.315 10.31 141.445 ;
		RECT	11.565 141.315 11.615 141.445 ;
		RECT	13.33 141.315 13.38 141.445 ;
		RECT	14.23 141.315 14.28 141.445 ;
		RECT	14.23 139.585 14.28 139.715 ;
		RECT	14.87 139.355 14.92 139.485 ;
		RECT	6.215 139.125 6.265 139.255 ;
		RECT	6.605 139.125 6.655 139.255 ;
		RECT	7.265 139.125 7.315 139.255 ;
		RECT	8.96 139.125 9.01 139.255 ;
		RECT	9.31 139.125 9.36 139.255 ;
		RECT	12.095 139.125 12.145 139.255 ;
		RECT	12.355 139.125 12.405 139.255 ;
		RECT	13.06 139.125 13.11 139.255 ;
		RECT	14.52 139.125 14.57 139.255 ;
		RECT	14.87 138.895 14.92 139.025 ;
		RECT	6.76 138.435 6.81 138.565 ;
		RECT	8.04 138.435 8.09 138.565 ;
		RECT	9.58 138.435 9.63 138.565 ;
		RECT	9.855 138.435 9.905 138.565 ;
		RECT	10.26 138.435 10.31 138.565 ;
		RECT	11.565 138.435 11.615 138.565 ;
		RECT	13.33 138.435 13.38 138.565 ;
		RECT	14.23 138.435 14.28 138.565 ;
		RECT	14.23 136.705 14.28 136.835 ;
		RECT	14.87 136.475 14.92 136.605 ;
		RECT	6.215 136.245 6.265 136.375 ;
		RECT	6.605 136.245 6.655 136.375 ;
		RECT	7.265 136.245 7.315 136.375 ;
		RECT	8.96 136.245 9.01 136.375 ;
		RECT	9.31 136.245 9.36 136.375 ;
		RECT	12.095 136.245 12.145 136.375 ;
		RECT	12.355 136.245 12.405 136.375 ;
		RECT	13.06 136.245 13.11 136.375 ;
		RECT	14.52 136.245 14.57 136.375 ;
		RECT	14.87 136.015 14.92 136.145 ;
		RECT	6.76 135.555 6.81 135.685 ;
		RECT	8.04 135.555 8.09 135.685 ;
		RECT	9.58 135.555 9.63 135.685 ;
		RECT	9.855 135.555 9.905 135.685 ;
		RECT	10.26 135.555 10.31 135.685 ;
		RECT	11.565 135.555 11.615 135.685 ;
		RECT	13.33 135.555 13.38 135.685 ;
		RECT	14.23 135.555 14.28 135.685 ;
		RECT	14.23 133.825 14.28 133.955 ;
		RECT	14.87 133.595 14.92 133.725 ;
		RECT	6.215 133.365 6.265 133.495 ;
		RECT	6.605 133.365 6.655 133.495 ;
		RECT	7.265 133.365 7.315 133.495 ;
		RECT	8.96 133.365 9.01 133.495 ;
		RECT	9.31 133.365 9.36 133.495 ;
		RECT	12.095 133.365 12.145 133.495 ;
		RECT	12.355 133.365 12.405 133.495 ;
		RECT	13.06 133.365 13.11 133.495 ;
		RECT	14.52 133.365 14.57 133.495 ;
		RECT	14.87 133.135 14.92 133.265 ;
		RECT	6.76 132.675 6.81 132.805 ;
		RECT	8.04 132.675 8.09 132.805 ;
		RECT	9.58 132.675 9.63 132.805 ;
		RECT	9.855 132.675 9.905 132.805 ;
		RECT	10.26 132.675 10.31 132.805 ;
		RECT	11.565 132.675 11.615 132.805 ;
		RECT	13.33 132.675 13.38 132.805 ;
		RECT	14.23 132.675 14.28 132.805 ;
		RECT	14.23 130.945 14.28 131.075 ;
		RECT	14.87 130.715 14.92 130.845 ;
		RECT	6.215 130.485 6.265 130.615 ;
		RECT	6.605 130.485 6.655 130.615 ;
		RECT	7.265 130.485 7.315 130.615 ;
		RECT	8.96 130.485 9.01 130.615 ;
		RECT	9.31 130.485 9.36 130.615 ;
		RECT	12.095 130.485 12.145 130.615 ;
		RECT	12.355 130.485 12.405 130.615 ;
		RECT	13.06 130.485 13.11 130.615 ;
		RECT	14.52 130.485 14.57 130.615 ;
		RECT	14.87 130.255 14.92 130.385 ;
		RECT	6.76 129.795 6.81 129.925 ;
		RECT	8.04 129.795 8.09 129.925 ;
		RECT	9.58 129.795 9.63 129.925 ;
		RECT	9.855 129.795 9.905 129.925 ;
		RECT	10.26 129.795 10.31 129.925 ;
		RECT	11.565 129.795 11.615 129.925 ;
		RECT	13.33 129.795 13.38 129.925 ;
		RECT	14.23 129.795 14.28 129.925 ;
		RECT	14.23 128.065 14.28 128.195 ;
		RECT	14.87 127.835 14.92 127.965 ;
		RECT	6.215 127.605 6.265 127.735 ;
		RECT	6.605 127.605 6.655 127.735 ;
		RECT	7.265 127.605 7.315 127.735 ;
		RECT	8.96 127.605 9.01 127.735 ;
		RECT	9.31 127.605 9.36 127.735 ;
		RECT	12.095 127.605 12.145 127.735 ;
		RECT	12.355 127.605 12.405 127.735 ;
		RECT	13.06 127.605 13.11 127.735 ;
		RECT	14.52 127.605 14.57 127.735 ;
		RECT	14.87 179.215 14.92 179.345 ;
		RECT	6.76 178.755 6.81 178.885 ;
		RECT	8.04 178.755 8.09 178.885 ;
		RECT	9.58 178.755 9.63 178.885 ;
		RECT	9.855 178.755 9.905 178.885 ;
		RECT	10.26 178.755 10.31 178.885 ;
		RECT	11.565 178.755 11.615 178.885 ;
		RECT	13.33 178.755 13.38 178.885 ;
		RECT	14.23 178.755 14.28 178.885 ;
		RECT	14.23 177.025 14.28 177.155 ;
		RECT	14.87 176.795 14.92 176.925 ;
		RECT	6.215 176.565 6.265 176.695 ;
		RECT	6.605 176.565 6.655 176.695 ;
		RECT	7.265 176.565 7.315 176.695 ;
		RECT	8.96 176.565 9.01 176.695 ;
		RECT	9.31 176.565 9.36 176.695 ;
		RECT	12.095 176.565 12.145 176.695 ;
		RECT	12.355 176.565 12.405 176.695 ;
		RECT	13.06 176.565 13.11 176.695 ;
		RECT	14.52 176.565 14.57 176.695 ;
		RECT	14.87 127.375 14.92 127.505 ;
		RECT	6.76 126.915 6.81 127.045 ;
		RECT	8.04 126.915 8.09 127.045 ;
		RECT	9.58 126.915 9.63 127.045 ;
		RECT	9.855 126.915 9.905 127.045 ;
		RECT	10.26 126.915 10.31 127.045 ;
		RECT	11.565 126.915 11.615 127.045 ;
		RECT	13.33 126.915 13.38 127.045 ;
		RECT	14.23 126.915 14.28 127.045 ;
		RECT	14.23 125.185 14.28 125.315 ;
		RECT	14.87 124.955 14.92 125.085 ;
		RECT	6.215 124.725 6.265 124.855 ;
		RECT	6.605 124.725 6.655 124.855 ;
		RECT	7.265 124.725 7.315 124.855 ;
		RECT	8.96 124.725 9.01 124.855 ;
		RECT	9.31 124.725 9.36 124.855 ;
		RECT	12.095 124.725 12.145 124.855 ;
		RECT	12.355 124.725 12.405 124.855 ;
		RECT	13.06 124.725 13.11 124.855 ;
		RECT	14.52 124.725 14.57 124.855 ;
		RECT	14.87 124.495 14.92 124.625 ;
		RECT	6.76 124.035 6.81 124.165 ;
		RECT	8.04 124.035 8.09 124.165 ;
		RECT	9.58 124.035 9.63 124.165 ;
		RECT	9.855 124.035 9.905 124.165 ;
		RECT	10.26 124.035 10.31 124.165 ;
		RECT	11.565 124.035 11.615 124.165 ;
		RECT	13.33 124.035 13.38 124.165 ;
		RECT	14.23 124.035 14.28 124.165 ;
		RECT	14.23 122.305 14.28 122.435 ;
		RECT	14.87 122.075 14.92 122.205 ;
		RECT	6.215 121.845 6.265 121.975 ;
		RECT	6.605 121.845 6.655 121.975 ;
		RECT	7.265 121.845 7.315 121.975 ;
		RECT	8.96 121.845 9.01 121.975 ;
		RECT	9.31 121.845 9.36 121.975 ;
		RECT	12.095 121.845 12.145 121.975 ;
		RECT	12.355 121.845 12.405 121.975 ;
		RECT	13.06 121.845 13.11 121.975 ;
		RECT	14.52 121.845 14.57 121.975 ;
		RECT	14.87 121.615 14.92 121.745 ;
		RECT	6.76 121.155 6.81 121.285 ;
		RECT	8.04 121.155 8.09 121.285 ;
		RECT	9.58 121.155 9.63 121.285 ;
		RECT	9.855 121.155 9.905 121.285 ;
		RECT	10.26 121.155 10.31 121.285 ;
		RECT	11.565 121.155 11.615 121.285 ;
		RECT	13.33 121.155 13.38 121.285 ;
		RECT	14.23 121.155 14.28 121.285 ;
		RECT	14.23 119.425 14.28 119.555 ;
		RECT	14.87 119.195 14.92 119.325 ;
		RECT	6.215 118.965 6.265 119.095 ;
		RECT	6.605 118.965 6.655 119.095 ;
		RECT	7.265 118.965 7.315 119.095 ;
		RECT	8.96 118.965 9.01 119.095 ;
		RECT	9.31 118.965 9.36 119.095 ;
		RECT	12.095 118.965 12.145 119.095 ;
		RECT	12.355 118.965 12.405 119.095 ;
		RECT	13.06 118.965 13.11 119.095 ;
		RECT	14.52 118.965 14.57 119.095 ;
		RECT	14.87 118.735 14.92 118.865 ;
		RECT	6.76 118.275 6.81 118.405 ;
		RECT	8.04 118.275 8.09 118.405 ;
		RECT	9.58 118.275 9.63 118.405 ;
		RECT	9.855 118.275 9.905 118.405 ;
		RECT	10.26 118.275 10.31 118.405 ;
		RECT	11.565 118.275 11.615 118.405 ;
		RECT	13.33 118.275 13.38 118.405 ;
		RECT	14.23 118.275 14.28 118.405 ;
		RECT	14.23 116.545 14.28 116.675 ;
		RECT	14.87 116.315 14.92 116.445 ;
		RECT	6.215 116.085 6.265 116.215 ;
		RECT	6.605 116.085 6.655 116.215 ;
		RECT	7.265 116.085 7.315 116.215 ;
		RECT	8.96 116.085 9.01 116.215 ;
		RECT	9.31 116.085 9.36 116.215 ;
		RECT	12.095 116.085 12.145 116.215 ;
		RECT	12.355 116.085 12.405 116.215 ;
		RECT	13.06 116.085 13.11 116.215 ;
		RECT	14.52 116.085 14.57 116.215 ;
		RECT	14.87 115.855 14.92 115.985 ;
		RECT	6.76 115.395 6.81 115.525 ;
		RECT	8.04 115.395 8.09 115.525 ;
		RECT	9.58 115.395 9.63 115.525 ;
		RECT	9.855 115.395 9.905 115.525 ;
		RECT	10.26 115.395 10.31 115.525 ;
		RECT	11.565 115.395 11.615 115.525 ;
		RECT	13.33 115.395 13.38 115.525 ;
		RECT	14.23 115.395 14.28 115.525 ;
		RECT	14.23 113.665 14.28 113.795 ;
		RECT	14.87 113.435 14.92 113.565 ;
		RECT	6.215 113.205 6.265 113.335 ;
		RECT	6.605 113.205 6.655 113.335 ;
		RECT	7.265 113.205 7.315 113.335 ;
		RECT	8.96 113.205 9.01 113.335 ;
		RECT	9.31 113.205 9.36 113.335 ;
		RECT	12.095 113.205 12.145 113.335 ;
		RECT	12.355 113.205 12.405 113.335 ;
		RECT	13.06 113.205 13.11 113.335 ;
		RECT	14.52 113.205 14.57 113.335 ;
		RECT	14.87 112.975 14.92 113.105 ;
		RECT	6.76 112.515 6.81 112.645 ;
		RECT	8.04 112.515 8.09 112.645 ;
		RECT	9.58 112.515 9.63 112.645 ;
		RECT	9.855 112.515 9.905 112.645 ;
		RECT	10.26 112.515 10.31 112.645 ;
		RECT	11.565 112.515 11.615 112.645 ;
		RECT	13.33 112.515 13.38 112.645 ;
		RECT	14.23 112.515 14.28 112.645 ;
		RECT	14.23 110.785 14.28 110.915 ;
		RECT	14.87 110.555 14.92 110.685 ;
		RECT	6.215 110.325 6.265 110.455 ;
		RECT	6.605 110.325 6.655 110.455 ;
		RECT	7.265 110.325 7.315 110.455 ;
		RECT	8.96 110.325 9.01 110.455 ;
		RECT	9.31 110.325 9.36 110.455 ;
		RECT	12.095 110.325 12.145 110.455 ;
		RECT	12.355 110.325 12.405 110.455 ;
		RECT	13.06 110.325 13.11 110.455 ;
		RECT	14.52 110.325 14.57 110.455 ;
		RECT	14.87 110.095 14.92 110.225 ;
		RECT	6.76 109.635 6.81 109.765 ;
		RECT	8.04 109.635 8.09 109.765 ;
		RECT	9.58 109.635 9.63 109.765 ;
		RECT	9.855 109.635 9.905 109.765 ;
		RECT	10.26 109.635 10.31 109.765 ;
		RECT	11.565 109.635 11.615 109.765 ;
		RECT	13.33 109.635 13.38 109.765 ;
		RECT	14.23 109.635 14.28 109.765 ;
		RECT	14.23 107.905 14.28 108.035 ;
		RECT	14.87 107.675 14.92 107.805 ;
		RECT	6.215 107.445 6.265 107.575 ;
		RECT	6.605 107.445 6.655 107.575 ;
		RECT	7.265 107.445 7.315 107.575 ;
		RECT	8.96 107.445 9.01 107.575 ;
		RECT	9.31 107.445 9.36 107.575 ;
		RECT	12.095 107.445 12.145 107.575 ;
		RECT	12.355 107.445 12.405 107.575 ;
		RECT	13.06 107.445 13.11 107.575 ;
		RECT	14.52 107.445 14.57 107.575 ;
		RECT	14.87 107.215 14.92 107.345 ;
		RECT	6.76 106.755 6.81 106.885 ;
		RECT	8.04 106.755 8.09 106.885 ;
		RECT	9.58 106.755 9.63 106.885 ;
		RECT	9.855 106.755 9.905 106.885 ;
		RECT	10.26 106.755 10.31 106.885 ;
		RECT	11.565 106.755 11.615 106.885 ;
		RECT	13.33 106.755 13.38 106.885 ;
		RECT	14.23 106.755 14.28 106.885 ;
		RECT	14.23 105.025 14.28 105.155 ;
		RECT	14.87 104.795 14.92 104.925 ;
		RECT	6.215 104.565 6.265 104.695 ;
		RECT	6.605 104.565 6.655 104.695 ;
		RECT	7.265 104.565 7.315 104.695 ;
		RECT	8.96 104.565 9.01 104.695 ;
		RECT	9.31 104.565 9.36 104.695 ;
		RECT	12.095 104.565 12.145 104.695 ;
		RECT	12.355 104.565 12.405 104.695 ;
		RECT	13.06 104.565 13.11 104.695 ;
		RECT	14.52 104.565 14.57 104.695 ;
		RECT	14.87 104.335 14.92 104.465 ;
		RECT	6.76 103.875 6.81 104.005 ;
		RECT	8.04 103.875 8.09 104.005 ;
		RECT	9.58 103.875 9.63 104.005 ;
		RECT	9.855 103.875 9.905 104.005 ;
		RECT	10.26 103.875 10.31 104.005 ;
		RECT	11.565 103.875 11.615 104.005 ;
		RECT	13.33 103.875 13.38 104.005 ;
		RECT	14.23 103.875 14.28 104.005 ;
		RECT	14.23 102.145 14.28 102.275 ;
		RECT	14.87 101.915 14.92 102.045 ;
		RECT	6.215 101.685 6.265 101.815 ;
		RECT	6.605 101.685 6.655 101.815 ;
		RECT	7.265 101.685 7.315 101.815 ;
		RECT	8.96 101.685 9.01 101.815 ;
		RECT	9.31 101.685 9.36 101.815 ;
		RECT	12.095 101.685 12.145 101.815 ;
		RECT	12.355 101.685 12.405 101.815 ;
		RECT	13.06 101.685 13.11 101.815 ;
		RECT	14.52 101.685 14.57 101.815 ;
		RECT	14.87 101.455 14.92 101.585 ;
		RECT	6.76 100.995 6.81 101.125 ;
		RECT	8.04 100.995 8.09 101.125 ;
		RECT	9.58 100.995 9.63 101.125 ;
		RECT	9.855 100.995 9.905 101.125 ;
		RECT	10.26 100.995 10.31 101.125 ;
		RECT	11.565 100.995 11.615 101.125 ;
		RECT	13.33 100.995 13.38 101.125 ;
		RECT	14.23 100.995 14.28 101.125 ;
		RECT	14.23 99.265 14.28 99.395 ;
		RECT	14.87 99.035 14.92 99.165 ;
		RECT	6.215 98.805 6.265 98.935 ;
		RECT	6.605 98.805 6.655 98.935 ;
		RECT	7.265 98.805 7.315 98.935 ;
		RECT	8.96 98.805 9.01 98.935 ;
		RECT	9.31 98.805 9.36 98.935 ;
		RECT	12.095 98.805 12.145 98.935 ;
		RECT	12.355 98.805 12.405 98.935 ;
		RECT	13.06 98.805 13.11 98.935 ;
		RECT	14.52 98.805 14.57 98.935 ;
		RECT	14.87 176.335 14.92 176.465 ;
		RECT	6.76 175.875 6.81 176.005 ;
		RECT	8.04 175.875 8.09 176.005 ;
		RECT	9.58 175.875 9.63 176.005 ;
		RECT	9.855 175.875 9.905 176.005 ;
		RECT	10.26 175.875 10.31 176.005 ;
		RECT	11.565 175.875 11.615 176.005 ;
		RECT	13.33 175.875 13.38 176.005 ;
		RECT	14.23 175.875 14.28 176.005 ;
		RECT	14.23 174.145 14.28 174.275 ;
		RECT	14.87 173.915 14.92 174.045 ;
		RECT	6.215 173.685 6.265 173.815 ;
		RECT	6.605 173.685 6.655 173.815 ;
		RECT	7.265 173.685 7.315 173.815 ;
		RECT	8.96 173.685 9.01 173.815 ;
		RECT	9.31 173.685 9.36 173.815 ;
		RECT	12.095 173.685 12.145 173.815 ;
		RECT	12.355 173.685 12.405 173.815 ;
		RECT	13.06 173.685 13.11 173.815 ;
		RECT	14.52 173.685 14.57 173.815 ;
		RECT	14.87 98.575 14.92 98.705 ;
		RECT	6.76 98.115 6.81 98.245 ;
		RECT	8.04 98.115 8.09 98.245 ;
		RECT	9.58 98.115 9.63 98.245 ;
		RECT	9.855 98.115 9.905 98.245 ;
		RECT	10.26 98.115 10.31 98.245 ;
		RECT	11.565 98.115 11.615 98.245 ;
		RECT	13.33 98.115 13.38 98.245 ;
		RECT	14.23 98.115 14.28 98.245 ;
		RECT	14.23 96.385 14.28 96.515 ;
		RECT	14.87 96.155 14.92 96.285 ;
		RECT	6.215 95.925 6.265 96.055 ;
		RECT	6.605 95.925 6.655 96.055 ;
		RECT	7.265 95.925 7.315 96.055 ;
		RECT	8.96 95.925 9.01 96.055 ;
		RECT	9.31 95.925 9.36 96.055 ;
		RECT	12.095 95.925 12.145 96.055 ;
		RECT	12.355 95.925 12.405 96.055 ;
		RECT	13.06 95.925 13.11 96.055 ;
		RECT	14.52 95.925 14.57 96.055 ;
		RECT	14.87 95.695 14.92 95.825 ;
		RECT	6.76 95.235 6.81 95.365 ;
		RECT	8.04 95.235 8.09 95.365 ;
		RECT	9.58 95.235 9.63 95.365 ;
		RECT	9.855 95.235 9.905 95.365 ;
		RECT	10.26 95.235 10.31 95.365 ;
		RECT	11.565 95.235 11.615 95.365 ;
		RECT	13.33 95.235 13.38 95.365 ;
		RECT	14.23 95.235 14.28 95.365 ;
		RECT	14.23 93.505 14.28 93.635 ;
		RECT	14.87 93.275 14.92 93.405 ;
		RECT	6.215 93.045 6.265 93.175 ;
		RECT	6.605 93.045 6.655 93.175 ;
		RECT	7.265 93.045 7.315 93.175 ;
		RECT	8.96 93.045 9.01 93.175 ;
		RECT	9.31 93.045 9.36 93.175 ;
		RECT	12.095 93.045 12.145 93.175 ;
		RECT	12.355 93.045 12.405 93.175 ;
		RECT	13.06 93.045 13.11 93.175 ;
		RECT	14.52 93.045 14.57 93.175 ;
		RECT	14.87 92.815 14.92 92.945 ;
		RECT	6.76 92.355 6.81 92.485 ;
		RECT	8.04 92.355 8.09 92.485 ;
		RECT	9.58 92.355 9.63 92.485 ;
		RECT	9.855 92.355 9.905 92.485 ;
		RECT	10.26 92.355 10.31 92.485 ;
		RECT	11.565 92.355 11.615 92.485 ;
		RECT	13.33 92.355 13.38 92.485 ;
		RECT	14.23 92.355 14.28 92.485 ;
		RECT	14.23 90.625 14.28 90.755 ;
		RECT	14.87 90.395 14.92 90.525 ;
		RECT	6.215 90.165 6.265 90.295 ;
		RECT	6.605 90.165 6.655 90.295 ;
		RECT	7.265 90.165 7.315 90.295 ;
		RECT	8.96 90.165 9.01 90.295 ;
		RECT	9.31 90.165 9.36 90.295 ;
		RECT	12.095 90.165 12.145 90.295 ;
		RECT	12.355 90.165 12.405 90.295 ;
		RECT	13.06 90.165 13.11 90.295 ;
		RECT	14.52 90.165 14.57 90.295 ;
		RECT	14.87 89.935 14.92 90.065 ;
		RECT	6.76 89.475 6.81 89.605 ;
		RECT	8.04 89.475 8.09 89.605 ;
		RECT	9.58 89.475 9.63 89.605 ;
		RECT	9.855 89.475 9.905 89.605 ;
		RECT	10.26 89.475 10.31 89.605 ;
		RECT	11.565 89.475 11.615 89.605 ;
		RECT	13.33 89.475 13.38 89.605 ;
		RECT	14.23 89.475 14.28 89.605 ;
		RECT	14.23 87.745 14.28 87.875 ;
		RECT	14.87 87.515 14.92 87.645 ;
		RECT	6.215 87.285 6.265 87.415 ;
		RECT	6.605 87.285 6.655 87.415 ;
		RECT	7.265 87.285 7.315 87.415 ;
		RECT	8.96 87.285 9.01 87.415 ;
		RECT	9.31 87.285 9.36 87.415 ;
		RECT	12.095 87.285 12.145 87.415 ;
		RECT	12.355 87.285 12.405 87.415 ;
		RECT	13.06 87.285 13.11 87.415 ;
		RECT	14.52 87.285 14.57 87.415 ;
		RECT	14.87 87.055 14.92 87.185 ;
		RECT	6.76 86.595 6.81 86.725 ;
		RECT	8.04 86.595 8.09 86.725 ;
		RECT	9.58 86.595 9.63 86.725 ;
		RECT	9.855 86.595 9.905 86.725 ;
		RECT	10.26 86.595 10.31 86.725 ;
		RECT	11.565 86.595 11.615 86.725 ;
		RECT	13.33 86.595 13.38 86.725 ;
		RECT	14.23 86.595 14.28 86.725 ;
		RECT	14.23 84.865 14.28 84.995 ;
		RECT	14.87 84.635 14.92 84.765 ;
		RECT	6.215 84.405 6.265 84.535 ;
		RECT	6.605 84.405 6.655 84.535 ;
		RECT	7.265 84.405 7.315 84.535 ;
		RECT	8.96 84.405 9.01 84.535 ;
		RECT	9.31 84.405 9.36 84.535 ;
		RECT	12.095 84.405 12.145 84.535 ;
		RECT	12.355 84.405 12.405 84.535 ;
		RECT	13.06 84.405 13.11 84.535 ;
		RECT	14.52 84.405 14.57 84.535 ;
		RECT	14.87 84.175 14.92 84.305 ;
		RECT	6.76 83.715 6.81 83.845 ;
		RECT	8.04 83.715 8.09 83.845 ;
		RECT	9.58 83.715 9.63 83.845 ;
		RECT	9.855 83.715 9.905 83.845 ;
		RECT	10.26 83.715 10.31 83.845 ;
		RECT	11.565 83.715 11.615 83.845 ;
		RECT	13.33 83.715 13.38 83.845 ;
		RECT	14.23 83.715 14.28 83.845 ;
		RECT	14.23 81.985 14.28 82.115 ;
		RECT	14.87 81.755 14.92 81.885 ;
		RECT	6.215 81.525 6.265 81.655 ;
		RECT	6.605 81.525 6.655 81.655 ;
		RECT	7.265 81.525 7.315 81.655 ;
		RECT	8.96 81.525 9.01 81.655 ;
		RECT	9.31 81.525 9.36 81.655 ;
		RECT	12.095 81.525 12.145 81.655 ;
		RECT	12.355 81.525 12.405 81.655 ;
		RECT	13.06 81.525 13.11 81.655 ;
		RECT	14.52 81.525 14.57 81.655 ;
		RECT	14.87 81.295 14.92 81.425 ;
		RECT	6.76 80.835 6.81 80.965 ;
		RECT	8.04 80.835 8.09 80.965 ;
		RECT	9.58 80.835 9.63 80.965 ;
		RECT	9.855 80.835 9.905 80.965 ;
		RECT	10.26 80.835 10.31 80.965 ;
		RECT	11.565 80.835 11.615 80.965 ;
		RECT	13.33 80.835 13.38 80.965 ;
		RECT	14.23 80.835 14.28 80.965 ;
		RECT	14.23 79.105 14.28 79.235 ;
		RECT	14.87 78.875 14.92 79.005 ;
		RECT	6.215 78.645 6.265 78.775 ;
		RECT	6.605 78.645 6.655 78.775 ;
		RECT	7.265 78.645 7.315 78.775 ;
		RECT	8.96 78.645 9.01 78.775 ;
		RECT	9.31 78.645 9.36 78.775 ;
		RECT	12.095 78.645 12.145 78.775 ;
		RECT	12.355 78.645 12.405 78.775 ;
		RECT	13.06 78.645 13.11 78.775 ;
		RECT	14.52 78.645 14.57 78.775 ;
		RECT	14.87 78.415 14.92 78.545 ;
		RECT	6.76 77.955 6.81 78.085 ;
		RECT	8.04 77.955 8.09 78.085 ;
		RECT	9.58 77.955 9.63 78.085 ;
		RECT	9.855 77.955 9.905 78.085 ;
		RECT	10.26 77.955 10.31 78.085 ;
		RECT	11.565 77.955 11.615 78.085 ;
		RECT	13.33 77.955 13.38 78.085 ;
		RECT	14.23 77.955 14.28 78.085 ;
		RECT	14.23 76.225 14.28 76.355 ;
		RECT	14.87 75.995 14.92 76.125 ;
		RECT	6.215 75.765 6.265 75.895 ;
		RECT	6.605 75.765 6.655 75.895 ;
		RECT	7.265 75.765 7.315 75.895 ;
		RECT	8.96 75.765 9.01 75.895 ;
		RECT	9.31 75.765 9.36 75.895 ;
		RECT	12.095 75.765 12.145 75.895 ;
		RECT	12.355 75.765 12.405 75.895 ;
		RECT	13.06 75.765 13.11 75.895 ;
		RECT	14.52 75.765 14.57 75.895 ;
		RECT	14.87 75.535 14.92 75.665 ;
		RECT	6.76 75.075 6.81 75.205 ;
		RECT	8.04 75.075 8.09 75.205 ;
		RECT	9.58 75.075 9.63 75.205 ;
		RECT	9.855 75.075 9.905 75.205 ;
		RECT	10.26 75.075 10.31 75.205 ;
		RECT	11.565 75.075 11.615 75.205 ;
		RECT	13.33 75.075 13.38 75.205 ;
		RECT	14.23 75.075 14.28 75.205 ;
		RECT	14.23 73.345 14.28 73.475 ;
		RECT	14.87 73.115 14.92 73.245 ;
		RECT	6.215 72.885 6.265 73.015 ;
		RECT	6.605 72.885 6.655 73.015 ;
		RECT	7.265 72.885 7.315 73.015 ;
		RECT	8.96 72.885 9.01 73.015 ;
		RECT	9.31 72.885 9.36 73.015 ;
		RECT	12.095 72.885 12.145 73.015 ;
		RECT	12.355 72.885 12.405 73.015 ;
		RECT	13.06 72.885 13.11 73.015 ;
		RECT	14.52 72.885 14.57 73.015 ;
		RECT	14.87 72.655 14.92 72.785 ;
		RECT	6.76 72.195 6.81 72.325 ;
		RECT	8.04 72.195 8.09 72.325 ;
		RECT	9.58 72.195 9.63 72.325 ;
		RECT	9.855 72.195 9.905 72.325 ;
		RECT	10.26 72.195 10.31 72.325 ;
		RECT	11.565 72.195 11.615 72.325 ;
		RECT	13.33 72.195 13.38 72.325 ;
		RECT	14.23 72.195 14.28 72.325 ;
		RECT	14.23 70.465 14.28 70.595 ;
		RECT	14.87 70.235 14.92 70.365 ;
		RECT	6.215 70.005 6.265 70.135 ;
		RECT	6.605 70.005 6.655 70.135 ;
		RECT	7.265 70.005 7.315 70.135 ;
		RECT	8.96 70.005 9.01 70.135 ;
		RECT	9.31 70.005 9.36 70.135 ;
		RECT	12.095 70.005 12.145 70.135 ;
		RECT	12.355 70.005 12.405 70.135 ;
		RECT	13.06 70.005 13.11 70.135 ;
		RECT	14.52 70.005 14.57 70.135 ;
		RECT	14.87 173.455 14.92 173.585 ;
		RECT	6.76 172.995 6.81 173.125 ;
		RECT	8.04 172.995 8.09 173.125 ;
		RECT	9.58 172.995 9.63 173.125 ;
		RECT	9.855 172.995 9.905 173.125 ;
		RECT	10.26 172.995 10.31 173.125 ;
		RECT	11.565 172.995 11.615 173.125 ;
		RECT	13.33 172.995 13.38 173.125 ;
		RECT	14.23 172.995 14.28 173.125 ;
		RECT	14.23 171.265 14.28 171.395 ;
		RECT	14.87 171.035 14.92 171.165 ;
		RECT	6.215 170.805 6.265 170.935 ;
		RECT	6.605 170.805 6.655 170.935 ;
		RECT	7.265 170.805 7.315 170.935 ;
		RECT	8.96 170.805 9.01 170.935 ;
		RECT	9.31 170.805 9.36 170.935 ;
		RECT	12.095 170.805 12.145 170.935 ;
		RECT	12.355 170.805 12.405 170.935 ;
		RECT	13.06 170.805 13.11 170.935 ;
		RECT	14.52 170.805 14.57 170.935 ;
		RECT	14.87 69.775 14.92 69.905 ;
		RECT	6.76 69.315 6.81 69.445 ;
		RECT	8.04 69.315 8.09 69.445 ;
		RECT	9.58 69.315 9.63 69.445 ;
		RECT	9.855 69.315 9.905 69.445 ;
		RECT	10.26 69.315 10.31 69.445 ;
		RECT	11.565 69.315 11.615 69.445 ;
		RECT	13.33 69.315 13.38 69.445 ;
		RECT	14.23 69.315 14.28 69.445 ;
		RECT	14.23 67.585 14.28 67.715 ;
		RECT	14.87 67.355 14.92 67.485 ;
		RECT	6.215 67.125 6.265 67.255 ;
		RECT	6.605 67.125 6.655 67.255 ;
		RECT	7.265 67.125 7.315 67.255 ;
		RECT	8.96 67.125 9.01 67.255 ;
		RECT	9.31 67.125 9.36 67.255 ;
		RECT	12.095 67.125 12.145 67.255 ;
		RECT	12.355 67.125 12.405 67.255 ;
		RECT	13.06 67.125 13.11 67.255 ;
		RECT	14.52 67.125 14.57 67.255 ;
		RECT	14.87 66.895 14.92 67.025 ;
		RECT	6.76 66.435 6.81 66.565 ;
		RECT	8.04 66.435 8.09 66.565 ;
		RECT	9.58 66.435 9.63 66.565 ;
		RECT	9.855 66.435 9.905 66.565 ;
		RECT	10.26 66.435 10.31 66.565 ;
		RECT	11.565 66.435 11.615 66.565 ;
		RECT	13.33 66.435 13.38 66.565 ;
		RECT	14.23 66.435 14.28 66.565 ;
		RECT	14.23 64.705 14.28 64.835 ;
		RECT	14.87 64.475 14.92 64.605 ;
		RECT	6.215 64.245 6.265 64.375 ;
		RECT	6.605 64.245 6.655 64.375 ;
		RECT	7.265 64.245 7.315 64.375 ;
		RECT	8.96 64.245 9.01 64.375 ;
		RECT	9.31 64.245 9.36 64.375 ;
		RECT	12.095 64.245 12.145 64.375 ;
		RECT	12.355 64.245 12.405 64.375 ;
		RECT	13.06 64.245 13.11 64.375 ;
		RECT	14.52 64.245 14.57 64.375 ;
		RECT	14.87 64.015 14.92 64.145 ;
		RECT	6.76 63.555 6.81 63.685 ;
		RECT	8.04 63.555 8.09 63.685 ;
		RECT	9.58 63.555 9.63 63.685 ;
		RECT	9.855 63.555 9.905 63.685 ;
		RECT	10.26 63.555 10.31 63.685 ;
		RECT	11.565 63.555 11.615 63.685 ;
		RECT	13.33 63.555 13.38 63.685 ;
		RECT	14.23 63.555 14.28 63.685 ;
		RECT	14.23 61.825 14.28 61.955 ;
		RECT	14.87 61.595 14.92 61.725 ;
		RECT	6.215 61.365 6.265 61.495 ;
		RECT	6.605 61.365 6.655 61.495 ;
		RECT	7.265 61.365 7.315 61.495 ;
		RECT	8.96 61.365 9.01 61.495 ;
		RECT	9.31 61.365 9.36 61.495 ;
		RECT	12.095 61.365 12.145 61.495 ;
		RECT	12.355 61.365 12.405 61.495 ;
		RECT	13.06 61.365 13.11 61.495 ;
		RECT	14.52 61.365 14.57 61.495 ;
		RECT	14.87 61.135 14.92 61.265 ;
		RECT	6.76 60.675 6.81 60.805 ;
		RECT	8.04 60.675 8.09 60.805 ;
		RECT	9.58 60.675 9.63 60.805 ;
		RECT	9.855 60.675 9.905 60.805 ;
		RECT	10.26 60.675 10.31 60.805 ;
		RECT	11.565 60.675 11.615 60.805 ;
		RECT	13.33 60.675 13.38 60.805 ;
		RECT	14.23 60.675 14.28 60.805 ;
		RECT	14.23 58.945 14.28 59.075 ;
		RECT	14.87 58.715 14.92 58.845 ;
		RECT	6.215 58.485 6.265 58.615 ;
		RECT	6.605 58.485 6.655 58.615 ;
		RECT	7.265 58.485 7.315 58.615 ;
		RECT	8.96 58.485 9.01 58.615 ;
		RECT	9.31 58.485 9.36 58.615 ;
		RECT	12.095 58.485 12.145 58.615 ;
		RECT	12.355 58.485 12.405 58.615 ;
		RECT	13.06 58.485 13.11 58.615 ;
		RECT	14.52 58.485 14.57 58.615 ;
		RECT	14.87 58.255 14.92 58.385 ;
		RECT	6.76 57.795 6.81 57.925 ;
		RECT	8.04 57.795 8.09 57.925 ;
		RECT	9.58 57.795 9.63 57.925 ;
		RECT	9.855 57.795 9.905 57.925 ;
		RECT	10.26 57.795 10.31 57.925 ;
		RECT	11.565 57.795 11.615 57.925 ;
		RECT	13.33 57.795 13.38 57.925 ;
		RECT	14.23 57.795 14.28 57.925 ;
		RECT	14.23 56.065 14.28 56.195 ;
		RECT	14.87 55.835 14.92 55.965 ;
		RECT	6.215 55.605 6.265 55.735 ;
		RECT	6.605 55.605 6.655 55.735 ;
		RECT	7.265 55.605 7.315 55.735 ;
		RECT	8.96 55.605 9.01 55.735 ;
		RECT	9.31 55.605 9.36 55.735 ;
		RECT	12.095 55.605 12.145 55.735 ;
		RECT	12.355 55.605 12.405 55.735 ;
		RECT	13.06 55.605 13.11 55.735 ;
		RECT	14.52 55.605 14.57 55.735 ;
		RECT	14.87 55.375 14.92 55.505 ;
		RECT	6.76 54.915 6.81 55.045 ;
		RECT	8.04 54.915 8.09 55.045 ;
		RECT	9.58 54.915 9.63 55.045 ;
		RECT	9.855 54.915 9.905 55.045 ;
		RECT	10.26 54.915 10.31 55.045 ;
		RECT	11.565 54.915 11.615 55.045 ;
		RECT	13.33 54.915 13.38 55.045 ;
		RECT	14.23 54.915 14.28 55.045 ;
		RECT	14.23 53.185 14.28 53.315 ;
		RECT	14.87 52.955 14.92 53.085 ;
		RECT	6.215 52.725 6.265 52.855 ;
		RECT	6.605 52.725 6.655 52.855 ;
		RECT	7.265 52.725 7.315 52.855 ;
		RECT	8.96 52.725 9.01 52.855 ;
		RECT	9.31 52.725 9.36 52.855 ;
		RECT	12.095 52.725 12.145 52.855 ;
		RECT	12.355 52.725 12.405 52.855 ;
		RECT	13.06 52.725 13.11 52.855 ;
		RECT	14.52 52.725 14.57 52.855 ;
		RECT	14.87 52.495 14.92 52.625 ;
		RECT	6.76 52.035 6.81 52.165 ;
		RECT	8.04 52.035 8.09 52.165 ;
		RECT	9.58 52.035 9.63 52.165 ;
		RECT	9.855 52.035 9.905 52.165 ;
		RECT	10.26 52.035 10.31 52.165 ;
		RECT	11.565 52.035 11.615 52.165 ;
		RECT	13.33 52.035 13.38 52.165 ;
		RECT	14.23 52.035 14.28 52.165 ;
		RECT	14.23 50.305 14.28 50.435 ;
		RECT	14.87 50.075 14.92 50.205 ;
		RECT	6.215 49.845 6.265 49.975 ;
		RECT	6.605 49.845 6.655 49.975 ;
		RECT	7.265 49.845 7.315 49.975 ;
		RECT	8.96 49.845 9.01 49.975 ;
		RECT	9.31 49.845 9.36 49.975 ;
		RECT	12.095 49.845 12.145 49.975 ;
		RECT	12.355 49.845 12.405 49.975 ;
		RECT	13.06 49.845 13.11 49.975 ;
		RECT	14.52 49.845 14.57 49.975 ;
		RECT	14.87 49.615 14.92 49.745 ;
		RECT	6.76 49.155 6.81 49.285 ;
		RECT	8.04 49.155 8.09 49.285 ;
		RECT	9.58 49.155 9.63 49.285 ;
		RECT	9.855 49.155 9.905 49.285 ;
		RECT	10.26 49.155 10.31 49.285 ;
		RECT	11.565 49.155 11.615 49.285 ;
		RECT	13.33 49.155 13.38 49.285 ;
		RECT	14.23 49.155 14.28 49.285 ;
		RECT	14.23 47.425 14.28 47.555 ;
		RECT	14.87 47.195 14.92 47.325 ;
		RECT	6.215 46.965 6.265 47.095 ;
		RECT	6.605 46.965 6.655 47.095 ;
		RECT	7.265 46.965 7.315 47.095 ;
		RECT	8.96 46.965 9.01 47.095 ;
		RECT	9.31 46.965 9.36 47.095 ;
		RECT	12.095 46.965 12.145 47.095 ;
		RECT	12.355 46.965 12.405 47.095 ;
		RECT	13.06 46.965 13.11 47.095 ;
		RECT	14.52 46.965 14.57 47.095 ;
		RECT	14.87 46.735 14.92 46.865 ;
		RECT	6.76 46.275 6.81 46.405 ;
		RECT	8.04 46.275 8.09 46.405 ;
		RECT	9.58 46.275 9.63 46.405 ;
		RECT	9.855 46.275 9.905 46.405 ;
		RECT	10.26 46.275 10.31 46.405 ;
		RECT	11.565 46.275 11.615 46.405 ;
		RECT	13.33 46.275 13.38 46.405 ;
		RECT	14.23 46.275 14.28 46.405 ;
		RECT	14.23 44.545 14.28 44.675 ;
		RECT	14.87 44.315 14.92 44.445 ;
		RECT	6.215 44.085 6.265 44.215 ;
		RECT	6.605 44.085 6.655 44.215 ;
		RECT	7.265 44.085 7.315 44.215 ;
		RECT	8.96 44.085 9.01 44.215 ;
		RECT	9.31 44.085 9.36 44.215 ;
		RECT	12.095 44.085 12.145 44.215 ;
		RECT	12.355 44.085 12.405 44.215 ;
		RECT	13.06 44.085 13.11 44.215 ;
		RECT	14.52 44.085 14.57 44.215 ;
		RECT	14.87 43.855 14.92 43.985 ;
		RECT	6.76 43.395 6.81 43.525 ;
		RECT	8.04 43.395 8.09 43.525 ;
		RECT	9.58 43.395 9.63 43.525 ;
		RECT	9.855 43.395 9.905 43.525 ;
		RECT	10.26 43.395 10.31 43.525 ;
		RECT	11.565 43.395 11.615 43.525 ;
		RECT	13.33 43.395 13.38 43.525 ;
		RECT	14.23 43.395 14.28 43.525 ;
		RECT	14.23 41.665 14.28 41.795 ;
		RECT	14.87 41.435 14.92 41.565 ;
		RECT	6.215 41.205 6.265 41.335 ;
		RECT	6.605 41.205 6.655 41.335 ;
		RECT	7.265 41.205 7.315 41.335 ;
		RECT	8.96 41.205 9.01 41.335 ;
		RECT	9.31 41.205 9.36 41.335 ;
		RECT	12.095 41.205 12.145 41.335 ;
		RECT	12.355 41.205 12.405 41.335 ;
		RECT	13.06 41.205 13.11 41.335 ;
		RECT	14.52 41.205 14.57 41.335 ;
		RECT	14.87 170.575 14.92 170.705 ;
		RECT	6.76 170.115 6.81 170.245 ;
		RECT	8.04 170.115 8.09 170.245 ;
		RECT	9.58 170.115 9.63 170.245 ;
		RECT	9.855 170.115 9.905 170.245 ;
		RECT	10.26 170.115 10.31 170.245 ;
		RECT	11.565 170.115 11.615 170.245 ;
		RECT	13.33 170.115 13.38 170.245 ;
		RECT	14.23 170.115 14.28 170.245 ;
		RECT	14.23 168.385 14.28 168.515 ;
		RECT	14.87 168.155 14.92 168.285 ;
		RECT	6.215 167.925 6.265 168.055 ;
		RECT	6.605 167.925 6.655 168.055 ;
		RECT	7.265 167.925 7.315 168.055 ;
		RECT	8.96 167.925 9.01 168.055 ;
		RECT	9.31 167.925 9.36 168.055 ;
		RECT	12.095 167.925 12.145 168.055 ;
		RECT	12.355 167.925 12.405 168.055 ;
		RECT	13.06 167.925 13.11 168.055 ;
		RECT	14.52 167.925 14.57 168.055 ;
		RECT	14.87 40.975 14.92 41.105 ;
		RECT	6.76 40.515 6.81 40.645 ;
		RECT	8.04 40.515 8.09 40.645 ;
		RECT	9.58 40.515 9.63 40.645 ;
		RECT	9.855 40.515 9.905 40.645 ;
		RECT	10.26 40.515 10.31 40.645 ;
		RECT	11.565 40.515 11.615 40.645 ;
		RECT	13.33 40.515 13.38 40.645 ;
		RECT	14.23 40.515 14.28 40.645 ;
		RECT	14.23 38.785 14.28 38.915 ;
		RECT	14.87 38.555 14.92 38.685 ;
		RECT	6.215 38.325 6.265 38.455 ;
		RECT	6.605 38.325 6.655 38.455 ;
		RECT	7.265 38.325 7.315 38.455 ;
		RECT	8.96 38.325 9.01 38.455 ;
		RECT	9.31 38.325 9.36 38.455 ;
		RECT	12.095 38.325 12.145 38.455 ;
		RECT	12.355 38.325 12.405 38.455 ;
		RECT	13.06 38.325 13.11 38.455 ;
		RECT	14.52 38.325 14.57 38.455 ;
		RECT	14.87 38.095 14.92 38.225 ;
		RECT	6.76 37.635 6.81 37.765 ;
		RECT	8.04 37.635 8.09 37.765 ;
		RECT	9.58 37.635 9.63 37.765 ;
		RECT	9.855 37.635 9.905 37.765 ;
		RECT	10.26 37.635 10.31 37.765 ;
		RECT	11.565 37.635 11.615 37.765 ;
		RECT	13.33 37.635 13.38 37.765 ;
		RECT	14.23 37.635 14.28 37.765 ;
		RECT	14.23 35.905 14.28 36.035 ;
		RECT	14.87 35.675 14.92 35.805 ;
		RECT	6.215 35.445 6.265 35.575 ;
		RECT	6.605 35.445 6.655 35.575 ;
		RECT	7.265 35.445 7.315 35.575 ;
		RECT	8.96 35.445 9.01 35.575 ;
		RECT	9.31 35.445 9.36 35.575 ;
		RECT	12.095 35.445 12.145 35.575 ;
		RECT	12.355 35.445 12.405 35.575 ;
		RECT	13.06 35.445 13.11 35.575 ;
		RECT	14.52 35.445 14.57 35.575 ;
		RECT	14.87 35.215 14.92 35.345 ;
		RECT	6.76 34.755 6.81 34.885 ;
		RECT	8.04 34.755 8.09 34.885 ;
		RECT	9.58 34.755 9.63 34.885 ;
		RECT	9.855 34.755 9.905 34.885 ;
		RECT	10.26 34.755 10.31 34.885 ;
		RECT	11.565 34.755 11.615 34.885 ;
		RECT	13.33 34.755 13.38 34.885 ;
		RECT	14.23 34.755 14.28 34.885 ;
		RECT	14.23 33.025 14.28 33.155 ;
		RECT	14.87 32.795 14.92 32.925 ;
		RECT	6.215 32.565 6.265 32.695 ;
		RECT	6.605 32.565 6.655 32.695 ;
		RECT	7.265 32.565 7.315 32.695 ;
		RECT	8.96 32.565 9.01 32.695 ;
		RECT	9.31 32.565 9.36 32.695 ;
		RECT	12.095 32.565 12.145 32.695 ;
		RECT	12.355 32.565 12.405 32.695 ;
		RECT	13.06 32.565 13.11 32.695 ;
		RECT	14.52 32.565 14.57 32.695 ;
		RECT	14.87 32.335 14.92 32.465 ;
		RECT	6.76 31.875 6.81 32.005 ;
		RECT	8.04 31.875 8.09 32.005 ;
		RECT	9.58 31.875 9.63 32.005 ;
		RECT	9.855 31.875 9.905 32.005 ;
		RECT	10.26 31.875 10.31 32.005 ;
		RECT	11.565 31.875 11.615 32.005 ;
		RECT	13.33 31.875 13.38 32.005 ;
		RECT	14.23 31.875 14.28 32.005 ;
		RECT	14.23 30.145 14.28 30.275 ;
		RECT	14.87 29.915 14.92 30.045 ;
		RECT	6.215 29.685 6.265 29.815 ;
		RECT	6.605 29.685 6.655 29.815 ;
		RECT	7.265 29.685 7.315 29.815 ;
		RECT	8.96 29.685 9.01 29.815 ;
		RECT	9.31 29.685 9.36 29.815 ;
		RECT	12.095 29.685 12.145 29.815 ;
		RECT	12.355 29.685 12.405 29.815 ;
		RECT	13.06 29.685 13.11 29.815 ;
		RECT	14.52 29.685 14.57 29.815 ;
		RECT	14.87 29.455 14.92 29.585 ;
		RECT	6.76 28.995 6.81 29.125 ;
		RECT	8.04 28.995 8.09 29.125 ;
		RECT	9.58 28.995 9.63 29.125 ;
		RECT	9.855 28.995 9.905 29.125 ;
		RECT	10.26 28.995 10.31 29.125 ;
		RECT	11.565 28.995 11.615 29.125 ;
		RECT	13.33 28.995 13.38 29.125 ;
		RECT	14.23 28.995 14.28 29.125 ;
		RECT	14.23 27.265 14.28 27.395 ;
		RECT	14.87 27.035 14.92 27.165 ;
		RECT	6.215 26.805 6.265 26.935 ;
		RECT	6.605 26.805 6.655 26.935 ;
		RECT	7.265 26.805 7.315 26.935 ;
		RECT	8.96 26.805 9.01 26.935 ;
		RECT	9.31 26.805 9.36 26.935 ;
		RECT	12.095 26.805 12.145 26.935 ;
		RECT	12.355 26.805 12.405 26.935 ;
		RECT	13.06 26.805 13.11 26.935 ;
		RECT	14.52 26.805 14.57 26.935 ;
		RECT	14.87 26.575 14.92 26.705 ;
		RECT	6.76 26.115 6.81 26.245 ;
		RECT	8.04 26.115 8.09 26.245 ;
		RECT	9.58 26.115 9.63 26.245 ;
		RECT	9.855 26.115 9.905 26.245 ;
		RECT	10.26 26.115 10.31 26.245 ;
		RECT	11.565 26.115 11.615 26.245 ;
		RECT	13.33 26.115 13.38 26.245 ;
		RECT	14.23 26.115 14.28 26.245 ;
		RECT	14.23 24.385 14.28 24.515 ;
		RECT	14.87 24.155 14.92 24.285 ;
		RECT	6.215 23.925 6.265 24.055 ;
		RECT	6.605 23.925 6.655 24.055 ;
		RECT	7.265 23.925 7.315 24.055 ;
		RECT	8.96 23.925 9.01 24.055 ;
		RECT	9.31 23.925 9.36 24.055 ;
		RECT	12.095 23.925 12.145 24.055 ;
		RECT	12.355 23.925 12.405 24.055 ;
		RECT	13.06 23.925 13.11 24.055 ;
		RECT	14.52 23.925 14.57 24.055 ;
		RECT	14.87 23.695 14.92 23.825 ;
		RECT	6.76 23.235 6.81 23.365 ;
		RECT	8.04 23.235 8.09 23.365 ;
		RECT	9.58 23.235 9.63 23.365 ;
		RECT	9.855 23.235 9.905 23.365 ;
		RECT	10.26 23.235 10.31 23.365 ;
		RECT	11.565 23.235 11.615 23.365 ;
		RECT	13.33 23.235 13.38 23.365 ;
		RECT	14.23 23.235 14.28 23.365 ;
		RECT	14.23 21.505 14.28 21.635 ;
		RECT	14.87 21.275 14.92 21.405 ;
		RECT	6.215 21.045 6.265 21.175 ;
		RECT	6.605 21.045 6.655 21.175 ;
		RECT	7.265 21.045 7.315 21.175 ;
		RECT	8.96 21.045 9.01 21.175 ;
		RECT	9.31 21.045 9.36 21.175 ;
		RECT	12.095 21.045 12.145 21.175 ;
		RECT	12.355 21.045 12.405 21.175 ;
		RECT	13.06 21.045 13.11 21.175 ;
		RECT	14.52 21.045 14.57 21.175 ;
		RECT	14.87 20.815 14.92 20.945 ;
		RECT	6.76 20.355 6.81 20.485 ;
		RECT	8.04 20.355 8.09 20.485 ;
		RECT	9.58 20.355 9.63 20.485 ;
		RECT	9.855 20.355 9.905 20.485 ;
		RECT	10.26 20.355 10.31 20.485 ;
		RECT	11.565 20.355 11.615 20.485 ;
		RECT	13.33 20.355 13.38 20.485 ;
		RECT	14.23 20.355 14.28 20.485 ;
		RECT	14.23 18.625 14.28 18.755 ;
		RECT	14.87 18.395 14.92 18.525 ;
		RECT	6.215 18.165 6.265 18.295 ;
		RECT	6.605 18.165 6.655 18.295 ;
		RECT	7.265 18.165 7.315 18.295 ;
		RECT	8.96 18.165 9.01 18.295 ;
		RECT	9.31 18.165 9.36 18.295 ;
		RECT	12.095 18.165 12.145 18.295 ;
		RECT	12.355 18.165 12.405 18.295 ;
		RECT	13.06 18.165 13.11 18.295 ;
		RECT	14.52 18.165 14.57 18.295 ;
		RECT	14.87 17.935 14.92 18.065 ;
		RECT	6.76 17.475 6.81 17.605 ;
		RECT	8.04 17.475 8.09 17.605 ;
		RECT	9.58 17.475 9.63 17.605 ;
		RECT	9.855 17.475 9.905 17.605 ;
		RECT	10.26 17.475 10.31 17.605 ;
		RECT	11.565 17.475 11.615 17.605 ;
		RECT	13.33 17.475 13.38 17.605 ;
		RECT	14.23 17.475 14.28 17.605 ;
		RECT	14.23 15.745 14.28 15.875 ;
		RECT	14.87 15.515 14.92 15.645 ;
		RECT	6.215 15.285 6.265 15.415 ;
		RECT	6.605 15.285 6.655 15.415 ;
		RECT	7.265 15.285 7.315 15.415 ;
		RECT	8.96 15.285 9.01 15.415 ;
		RECT	9.31 15.285 9.36 15.415 ;
		RECT	12.095 15.285 12.145 15.415 ;
		RECT	12.355 15.285 12.405 15.415 ;
		RECT	13.06 15.285 13.11 15.415 ;
		RECT	14.52 15.285 14.57 15.415 ;
		RECT	14.87 15.055 14.92 15.185 ;
		RECT	6.76 14.595 6.81 14.725 ;
		RECT	8.04 14.595 8.09 14.725 ;
		RECT	9.58 14.595 9.63 14.725 ;
		RECT	9.855 14.595 9.905 14.725 ;
		RECT	10.26 14.595 10.31 14.725 ;
		RECT	11.565 14.595 11.615 14.725 ;
		RECT	13.33 14.595 13.38 14.725 ;
		RECT	14.23 14.595 14.28 14.725 ;
		RECT	14.23 12.865 14.28 12.995 ;
		RECT	14.87 12.635 14.92 12.765 ;
		RECT	6.215 12.405 6.265 12.535 ;
		RECT	6.605 12.405 6.655 12.535 ;
		RECT	7.265 12.405 7.315 12.535 ;
		RECT	8.96 12.405 9.01 12.535 ;
		RECT	9.31 12.405 9.36 12.535 ;
		RECT	12.095 12.405 12.145 12.535 ;
		RECT	12.355 12.405 12.405 12.535 ;
		RECT	13.06 12.405 13.11 12.535 ;
		RECT	14.52 12.405 14.57 12.535 ;
		RECT	14.87 167.695 14.92 167.825 ;
		RECT	6.76 167.235 6.81 167.365 ;
		RECT	8.04 167.235 8.09 167.365 ;
		RECT	9.58 167.235 9.63 167.365 ;
		RECT	9.855 167.235 9.905 167.365 ;
		RECT	10.26 167.235 10.31 167.365 ;
		RECT	11.565 167.235 11.615 167.365 ;
		RECT	13.33 167.235 13.38 167.365 ;
		RECT	14.23 167.235 14.28 167.365 ;
		RECT	14.23 165.505 14.28 165.635 ;
		RECT	14.87 165.275 14.92 165.405 ;
		RECT	6.215 165.045 6.265 165.175 ;
		RECT	6.605 165.045 6.655 165.175 ;
		RECT	7.265 165.045 7.315 165.175 ;
		RECT	8.96 165.045 9.01 165.175 ;
		RECT	9.31 165.045 9.36 165.175 ;
		RECT	12.095 165.045 12.145 165.175 ;
		RECT	12.355 165.045 12.405 165.175 ;
		RECT	13.06 165.045 13.11 165.175 ;
		RECT	14.52 165.045 14.57 165.175 ;
		RECT	14.87 12.175 14.92 12.305 ;
		RECT	6.76 11.715 6.81 11.845 ;
		RECT	8.04 11.715 8.09 11.845 ;
		RECT	9.58 11.715 9.63 11.845 ;
		RECT	9.855 11.715 9.905 11.845 ;
		RECT	10.26 11.715 10.31 11.845 ;
		RECT	11.565 11.715 11.615 11.845 ;
		RECT	13.33 11.715 13.38 11.845 ;
		RECT	14.23 11.715 14.28 11.845 ;
		RECT	14.23 9.985 14.28 10.115 ;
		RECT	14.87 9.755 14.92 9.885 ;
		RECT	6.215 9.525 6.265 9.655 ;
		RECT	6.605 9.525 6.655 9.655 ;
		RECT	7.265 9.525 7.315 9.655 ;
		RECT	8.96 9.525 9.01 9.655 ;
		RECT	9.31 9.525 9.36 9.655 ;
		RECT	12.095 9.525 12.145 9.655 ;
		RECT	12.355 9.525 12.405 9.655 ;
		RECT	13.06 9.525 13.11 9.655 ;
		RECT	14.52 9.525 14.57 9.655 ;
		RECT	14.87 9.295 14.92 9.425 ;
		RECT	6.76 8.835 6.81 8.965 ;
		RECT	8.04 8.835 8.09 8.965 ;
		RECT	9.58 8.835 9.63 8.965 ;
		RECT	9.855 8.835 9.905 8.965 ;
		RECT	10.26 8.835 10.31 8.965 ;
		RECT	11.565 8.835 11.615 8.965 ;
		RECT	13.33 8.835 13.38 8.965 ;
		RECT	14.23 8.835 14.28 8.965 ;
		RECT	14.23 7.105 14.28 7.235 ;
		RECT	14.87 6.875 14.92 7.005 ;
		RECT	6.215 6.645 6.265 6.775 ;
		RECT	6.605 6.645 6.655 6.775 ;
		RECT	7.265 6.645 7.315 6.775 ;
		RECT	8.96 6.645 9.01 6.775 ;
		RECT	9.31 6.645 9.36 6.775 ;
		RECT	12.095 6.645 12.145 6.775 ;
		RECT	12.355 6.645 12.405 6.775 ;
		RECT	13.06 6.645 13.11 6.775 ;
		RECT	14.52 6.645 14.57 6.775 ;
		RECT	14.87 6.415 14.92 6.545 ;
		RECT	6.76 5.955 6.81 6.085 ;
		RECT	8.04 5.955 8.09 6.085 ;
		RECT	9.58 5.955 9.63 6.085 ;
		RECT	9.855 5.955 9.905 6.085 ;
		RECT	10.26 5.955 10.31 6.085 ;
		RECT	11.565 5.955 11.615 6.085 ;
		RECT	13.33 5.955 13.38 6.085 ;
		RECT	14.23 5.955 14.28 6.085 ;
		RECT	14.23 4.225 14.28 4.355 ;
		RECT	14.87 3.995 14.92 4.125 ;
		RECT	6.215 3.765 6.265 3.895 ;
		RECT	6.605 3.765 6.655 3.895 ;
		RECT	7.265 3.765 7.315 3.895 ;
		RECT	8.96 3.765 9.01 3.895 ;
		RECT	9.31 3.765 9.36 3.895 ;
		RECT	12.095 3.765 12.145 3.895 ;
		RECT	12.355 3.765 12.405 3.895 ;
		RECT	13.06 3.765 13.11 3.895 ;
		RECT	14.52 3.765 14.57 3.895 ;
		RECT	14.87 164.815 14.92 164.945 ;
		RECT	6.76 164.355 6.81 164.485 ;
		RECT	8.04 164.355 8.09 164.485 ;
		RECT	9.58 164.355 9.63 164.485 ;
		RECT	9.855 164.355 9.905 164.485 ;
		RECT	10.26 164.355 10.31 164.485 ;
		RECT	11.565 164.355 11.615 164.485 ;
		RECT	13.33 164.355 13.38 164.485 ;
		RECT	14.23 164.355 14.28 164.485 ;
		RECT	14.23 162.625 14.28 162.755 ;
		RECT	14.87 162.395 14.92 162.525 ;
		RECT	6.215 162.165 6.265 162.295 ;
		RECT	6.605 162.165 6.655 162.295 ;
		RECT	7.265 162.165 7.315 162.295 ;
		RECT	8.96 162.165 9.01 162.295 ;
		RECT	9.31 162.165 9.36 162.295 ;
		RECT	12.095 162.165 12.145 162.295 ;
		RECT	12.355 162.165 12.405 162.295 ;
		RECT	13.06 162.165 13.11 162.295 ;
		RECT	14.52 162.165 14.57 162.295 ;
		RECT	14.87 161.935 14.92 162.065 ;
		RECT	6.76 161.475 6.81 161.605 ;
		RECT	8.04 161.475 8.09 161.605 ;
		RECT	9.58 161.475 9.63 161.605 ;
		RECT	9.855 161.475 9.905 161.605 ;
		RECT	10.26 161.475 10.31 161.605 ;
		RECT	11.565 161.475 11.615 161.605 ;
		RECT	13.33 161.475 13.38 161.605 ;
		RECT	14.23 161.475 14.28 161.605 ;
		RECT	14.23 159.745 14.28 159.875 ;
		RECT	14.87 159.515 14.92 159.645 ;
		RECT	6.215 159.285 6.265 159.415 ;
		RECT	6.605 159.285 6.655 159.415 ;
		RECT	7.265 159.285 7.315 159.415 ;
		RECT	8.96 159.285 9.01 159.415 ;
		RECT	9.31 159.285 9.36 159.415 ;
		RECT	12.095 159.285 12.145 159.415 ;
		RECT	12.355 159.285 12.405 159.415 ;
		RECT	13.06 159.285 13.11 159.415 ;
		RECT	14.52 159.285 14.57 159.415 ;
		RECT	14.87 159.055 14.92 159.185 ;
		RECT	6.76 158.595 6.81 158.725 ;
		RECT	8.04 158.595 8.09 158.725 ;
		RECT	9.58 158.595 9.63 158.725 ;
		RECT	9.855 158.595 9.905 158.725 ;
		RECT	10.26 158.595 10.31 158.725 ;
		RECT	11.565 158.595 11.615 158.725 ;
		RECT	13.33 158.595 13.38 158.725 ;
		RECT	14.23 158.595 14.28 158.725 ;
		RECT	14.23 156.865 14.28 156.995 ;
		RECT	14.87 156.635 14.92 156.765 ;
		RECT	6.215 156.405 6.265 156.535 ;
		RECT	6.605 156.405 6.655 156.535 ;
		RECT	7.265 156.405 7.315 156.535 ;
		RECT	8.96 156.405 9.01 156.535 ;
		RECT	9.31 156.405 9.36 156.535 ;
		RECT	12.095 156.405 12.145 156.535 ;
		RECT	12.355 156.405 12.405 156.535 ;
		RECT	13.06 156.405 13.11 156.535 ;
		RECT	14.52 156.405 14.57 156.535 ;
		RECT	14.87 3.535 14.92 3.665 ;
		RECT	6.76 3.075 6.81 3.205 ;
		RECT	8.04 3.075 8.09 3.205 ;
		RECT	9.58 3.075 9.63 3.205 ;
		RECT	9.855 3.075 9.905 3.205 ;
		RECT	10.26 3.075 10.31 3.205 ;
		RECT	11.565 3.075 11.615 3.205 ;
		RECT	13.33 3.075 13.38 3.205 ;
		RECT	14.23 3.075 14.28 3.205 ;
		RECT	14.23 1.345 14.28 1.475 ;
		RECT	14.87 1.115 14.92 1.245 ;
		RECT	6.215 0.885 6.265 1.015 ;
		RECT	6.605 0.885 6.655 1.015 ;
		RECT	7.265 0.885 7.315 1.015 ;
		RECT	8.96 0.885 9.01 1.015 ;
		RECT	9.31 0.885 9.36 1.015 ;
		RECT	12.095 0.885 12.145 1.015 ;
		RECT	12.355 0.885 12.405 1.015 ;
		RECT	13.06 0.885 13.11 1.015 ;
		RECT	14.52 0.885 14.57 1.015 ;
		RECT	14.87 184.975 14.92 185.105 ;
		RECT	6.76 184.515 6.81 184.645 ;
		RECT	8.04 184.515 8.09 184.645 ;
		RECT	9.58 184.515 9.63 184.645 ;
		RECT	9.855 184.515 9.905 184.645 ;
		RECT	10.26 184.515 10.31 184.645 ;
		RECT	11.565 184.515 11.615 184.645 ;
		RECT	13.33 184.515 13.38 184.645 ;
		RECT	14.23 184.515 14.28 184.645 ;
		RECT	14.23 182.785 14.28 182.915 ;
		RECT	14.87 182.555 14.92 182.685 ;
		RECT	6.215 182.325 6.265 182.455 ;
		RECT	6.605 182.325 6.655 182.455 ;
		RECT	7.265 182.325 7.315 182.455 ;
		RECT	8.96 182.325 9.01 182.455 ;
		RECT	9.31 182.325 9.36 182.455 ;
		RECT	12.095 182.325 12.145 182.455 ;
		RECT	12.355 182.325 12.405 182.455 ;
		RECT	13.06 182.325 13.11 182.455 ;
		RECT	14.52 182.325 14.57 182.455 ;
		RECT	4.38 0.195 4.43 0.325 ;
		RECT	6.175 0.195 6.225 0.325 ;
		RECT	14.52 0.195 14.57 0.325 ;
		RECT	3.6 0.655 3.65 0.785 ;
		RECT	1.44 0.195 1.49 0.325 ;
		RECT	2.11 0.195 2.16 0.325 ;
		RECT	3.09 0.195 3.14 0.325 ;
		RECT	7.73 0.195 7.78 0.325 ;
		RECT	14.68 0.195 14.73 0.325 ;
		RECT	14.34 0.425 14.39 0.555 ;
		RECT	9.1 0.655 9.15 0.785 ;
		RECT	10.81 0.655 10.86 0.785 ;
		RECT	0.435 0.655 0.485 0.785 ;
		RECT	0.62 0.195 0.67 0.325 ;
		RECT	4.19 0.195 4.24 0.325 ;
		RECT	2.72 0.655 2.77 0.785 ;
		RECT	0.9 179.445 0.95 179.575 ;
		RECT	0.9 153.525 0.95 153.655 ;
		RECT	0.9 150.645 0.95 150.775 ;
		RECT	0.9 147.765 0.95 147.895 ;
		RECT	0.9 144.885 0.95 145.015 ;
		RECT	0.9 142.005 0.95 142.135 ;
		RECT	0.9 139.125 0.95 139.255 ;
		RECT	0.9 136.245 0.95 136.375 ;
		RECT	0.9 133.365 0.95 133.495 ;
		RECT	0.9 130.485 0.95 130.615 ;
		RECT	0.9 127.605 0.95 127.735 ;
		RECT	0.9 176.565 0.95 176.695 ;
		RECT	0.9 124.725 0.95 124.855 ;
		RECT	0.9 121.845 0.95 121.975 ;
		RECT	0.9 118.965 0.95 119.095 ;
		RECT	0.9 116.085 0.95 116.215 ;
		RECT	0.9 113.205 0.95 113.335 ;
		RECT	0.9 110.325 0.95 110.455 ;
		RECT	0.9 107.445 0.95 107.575 ;
		RECT	0.9 104.565 0.95 104.695 ;
		RECT	0.9 101.685 0.95 101.815 ;
		RECT	0.9 98.805 0.95 98.935 ;
		RECT	0.9 173.685 0.95 173.815 ;
		RECT	0.9 95.925 0.95 96.055 ;
		RECT	0.9 93.045 0.95 93.175 ;
		RECT	0.9 90.165 0.95 90.295 ;
		RECT	0.9 87.285 0.95 87.415 ;
		RECT	0.9 84.405 0.95 84.535 ;
		RECT	0.9 81.525 0.95 81.655 ;
		RECT	0.9 78.645 0.95 78.775 ;
		RECT	0.9 75.765 0.95 75.895 ;
		RECT	0.9 72.885 0.95 73.015 ;
		RECT	0.9 70.005 0.95 70.135 ;
		RECT	0.9 170.805 0.95 170.935 ;
		RECT	0.9 67.125 0.95 67.255 ;
		RECT	0.9 64.245 0.95 64.375 ;
		RECT	0.9 61.365 0.95 61.495 ;
		RECT	0.9 58.485 0.95 58.615 ;
		RECT	0.9 55.605 0.95 55.735 ;
		RECT	0.9 52.725 0.95 52.855 ;
		RECT	0.9 49.845 0.95 49.975 ;
		RECT	0.9 46.965 0.95 47.095 ;
		RECT	0.9 44.085 0.95 44.215 ;
		RECT	0.9 41.205 0.95 41.335 ;
		RECT	0.9 167.925 0.95 168.055 ;
		RECT	0.9 38.325 0.95 38.455 ;
		RECT	0.9 35.445 0.95 35.575 ;
		RECT	0.9 32.565 0.95 32.695 ;
		RECT	0.9 29.685 0.95 29.815 ;
		RECT	0.9 26.805 0.95 26.935 ;
		RECT	0.9 23.925 0.95 24.055 ;
		RECT	0.9 21.045 0.95 21.175 ;
		RECT	0.9 18.165 0.95 18.295 ;
		RECT	0.9 15.285 0.95 15.415 ;
		RECT	0.9 12.405 0.95 12.535 ;
		RECT	0.9 165.045 0.95 165.175 ;
		RECT	0.9 9.525 0.95 9.655 ;
		RECT	0.9 6.645 0.95 6.775 ;
		RECT	0.9 3.765 0.95 3.895 ;
		RECT	0.9 162.165 0.95 162.295 ;
		RECT	0.9 159.285 0.95 159.415 ;
		RECT	0.9 156.405 0.95 156.535 ;
		RECT	0.9 0.885 0.95 1.015 ;
		RECT	0.9 182.325 0.95 182.455 ;
		RECT	2.72 184.975 2.77 185.105 ;
		RECT	2.72 182.555 2.77 182.685 ;
		RECT	2.72 156.175 2.77 156.305 ;
		RECT	2.72 153.755 2.77 153.885 ;
		RECT	2.72 153.295 2.77 153.425 ;
		RECT	2.72 150.875 2.77 151.005 ;
		RECT	2.72 150.415 2.77 150.545 ;
		RECT	2.72 147.995 2.77 148.125 ;
		RECT	2.72 147.535 2.77 147.665 ;
		RECT	2.72 145.115 2.77 145.245 ;
		RECT	2.72 144.655 2.77 144.785 ;
		RECT	2.72 142.235 2.77 142.365 ;
		RECT	2.72 141.775 2.77 141.905 ;
		RECT	2.72 139.355 2.77 139.485 ;
		RECT	2.72 138.895 2.77 139.025 ;
		RECT	2.72 136.475 2.77 136.605 ;
		RECT	2.72 136.015 2.77 136.145 ;
		RECT	2.72 133.595 2.77 133.725 ;
		RECT	2.72 133.135 2.77 133.265 ;
		RECT	2.72 130.715 2.77 130.845 ;
		RECT	2.72 130.255 2.77 130.385 ;
		RECT	2.72 127.835 2.77 127.965 ;
		RECT	2.72 182.095 2.77 182.225 ;
		RECT	2.72 179.675 2.77 179.805 ;
		RECT	2.72 127.375 2.77 127.505 ;
		RECT	2.72 124.955 2.77 125.085 ;
		RECT	2.72 124.495 2.77 124.625 ;
		RECT	2.72 122.075 2.77 122.205 ;
		RECT	2.72 121.615 2.77 121.745 ;
		RECT	2.72 119.195 2.77 119.325 ;
		RECT	2.72 118.735 2.77 118.865 ;
		RECT	2.72 116.315 2.77 116.445 ;
		RECT	2.72 115.855 2.77 115.985 ;
		RECT	2.72 113.435 2.77 113.565 ;
		RECT	2.72 112.975 2.77 113.105 ;
		RECT	2.72 110.555 2.77 110.685 ;
		RECT	2.72 110.095 2.77 110.225 ;
		RECT	2.72 107.675 2.77 107.805 ;
		RECT	2.72 107.215 2.77 107.345 ;
		RECT	2.72 104.795 2.77 104.925 ;
		RECT	2.72 104.335 2.77 104.465 ;
		RECT	2.72 101.915 2.77 102.045 ;
		RECT	2.72 101.455 2.77 101.585 ;
		RECT	2.72 99.035 2.77 99.165 ;
		RECT	2.72 179.215 2.77 179.345 ;
		RECT	2.72 176.795 2.77 176.925 ;
		RECT	2.72 98.575 2.77 98.705 ;
		RECT	2.72 96.155 2.77 96.285 ;
		RECT	2.72 95.695 2.77 95.825 ;
		RECT	2.72 93.275 2.77 93.405 ;
		RECT	2.72 92.815 2.77 92.945 ;
		RECT	2.72 90.395 2.77 90.525 ;
		RECT	2.72 89.935 2.77 90.065 ;
		RECT	2.72 87.515 2.77 87.645 ;
		RECT	2.72 87.055 2.77 87.185 ;
		RECT	2.72 84.635 2.77 84.765 ;
		RECT	2.72 84.175 2.77 84.305 ;
		RECT	2.72 81.755 2.77 81.885 ;
		RECT	2.72 81.295 2.77 81.425 ;
		RECT	2.72 78.875 2.77 79.005 ;
		RECT	2.72 78.415 2.77 78.545 ;
		RECT	2.72 75.995 2.77 76.125 ;
		RECT	2.72 75.535 2.77 75.665 ;
		RECT	2.72 73.115 2.77 73.245 ;
		RECT	2.72 72.655 2.77 72.785 ;
		RECT	2.72 70.235 2.77 70.365 ;
		RECT	2.72 176.335 2.77 176.465 ;
		RECT	2.72 173.915 2.77 174.045 ;
		RECT	2.72 69.775 2.77 69.905 ;
		RECT	2.72 67.355 2.77 67.485 ;
		RECT	2.72 66.895 2.77 67.025 ;
		RECT	2.72 64.475 2.77 64.605 ;
		RECT	2.72 64.015 2.77 64.145 ;
		RECT	2.72 61.595 2.77 61.725 ;
		RECT	2.72 61.135 2.77 61.265 ;
		RECT	2.72 58.715 2.77 58.845 ;
		RECT	2.72 58.255 2.77 58.385 ;
		RECT	2.72 55.835 2.77 55.965 ;
		RECT	2.72 55.375 2.77 55.505 ;
		RECT	2.72 52.955 2.77 53.085 ;
		RECT	2.72 52.495 2.77 52.625 ;
		RECT	2.72 50.075 2.77 50.205 ;
		RECT	2.72 49.615 2.77 49.745 ;
		RECT	2.72 47.195 2.77 47.325 ;
		RECT	2.72 46.735 2.77 46.865 ;
		RECT	2.72 44.315 2.77 44.445 ;
		RECT	2.72 43.855 2.77 43.985 ;
		RECT	2.72 41.435 2.77 41.565 ;
		RECT	2.72 173.455 2.77 173.585 ;
		RECT	2.72 171.035 2.77 171.165 ;
		RECT	2.72 40.975 2.77 41.105 ;
		RECT	2.72 38.555 2.77 38.685 ;
		RECT	2.72 38.095 2.77 38.225 ;
		RECT	2.72 35.675 2.77 35.805 ;
		RECT	2.72 35.215 2.77 35.345 ;
		RECT	2.72 32.795 2.77 32.925 ;
		RECT	2.72 32.335 2.77 32.465 ;
		RECT	2.72 29.915 2.77 30.045 ;
		RECT	2.72 29.455 2.77 29.585 ;
		RECT	2.72 27.035 2.77 27.165 ;
		RECT	2.72 26.575 2.77 26.705 ;
		RECT	2.72 24.155 2.77 24.285 ;
		RECT	2.72 23.695 2.77 23.825 ;
		RECT	2.72 21.275 2.77 21.405 ;
		RECT	2.72 20.815 2.77 20.945 ;
		RECT	2.72 18.395 2.77 18.525 ;
		RECT	2.72 17.935 2.77 18.065 ;
		RECT	2.72 15.515 2.77 15.645 ;
		RECT	2.72 15.055 2.77 15.185 ;
		RECT	2.72 12.635 2.77 12.765 ;
		RECT	2.72 170.575 2.77 170.705 ;
		RECT	2.72 168.155 2.77 168.285 ;
		RECT	2.72 12.175 2.77 12.305 ;
		RECT	2.72 9.755 2.77 9.885 ;
		RECT	2.72 9.295 2.77 9.425 ;
		RECT	2.72 6.875 2.77 7.005 ;
		RECT	2.72 6.415 2.77 6.545 ;
		RECT	2.72 3.995 2.77 4.125 ;
		RECT	2.72 3.535 2.77 3.665 ;
		RECT	2.72 1.115 2.77 1.245 ;
		RECT	2.72 167.695 2.77 167.825 ;
		RECT	2.72 165.275 2.77 165.405 ;
		RECT	2.72 164.815 2.77 164.945 ;
		RECT	2.72 162.395 2.77 162.525 ;
		RECT	2.72 161.935 2.77 162.065 ;
		RECT	2.72 159.515 2.77 159.645 ;
		RECT	2.72 159.055 2.77 159.185 ;
		RECT	2.72 156.635 2.77 156.765 ;
		RECT	1.625 184.975 1.675 185.105 ;
		RECT	1.92 184.975 1.97 185.105 ;
		RECT	5.05 184.975 5.1 185.105 ;
		RECT	3.6 184.515 3.65 184.645 ;
		RECT	1.625 182.555 1.675 182.685 ;
		RECT	1.92 182.555 1.97 182.685 ;
		RECT	5.05 182.555 5.1 182.685 ;
		RECT	1.625 156.175 1.675 156.305 ;
		RECT	1.92 156.175 1.97 156.305 ;
		RECT	5.05 156.175 5.1 156.305 ;
		RECT	3.6 155.715 3.65 155.845 ;
		RECT	1.625 153.755 1.675 153.885 ;
		RECT	1.92 153.755 1.97 153.885 ;
		RECT	5.05 153.755 5.1 153.885 ;
		RECT	1.625 153.295 1.675 153.425 ;
		RECT	1.92 153.295 1.97 153.425 ;
		RECT	5.05 153.295 5.1 153.425 ;
		RECT	3.6 152.835 3.65 152.965 ;
		RECT	1.625 150.875 1.675 151.005 ;
		RECT	1.92 150.875 1.97 151.005 ;
		RECT	5.05 150.875 5.1 151.005 ;
		RECT	1.625 150.415 1.675 150.545 ;
		RECT	1.92 150.415 1.97 150.545 ;
		RECT	5.05 150.415 5.1 150.545 ;
		RECT	3.6 149.955 3.65 150.085 ;
		RECT	1.625 147.995 1.675 148.125 ;
		RECT	1.92 147.995 1.97 148.125 ;
		RECT	5.05 147.995 5.1 148.125 ;
		RECT	1.625 147.535 1.675 147.665 ;
		RECT	1.92 147.535 1.97 147.665 ;
		RECT	5.05 147.535 5.1 147.665 ;
		RECT	3.6 147.075 3.65 147.205 ;
		RECT	1.625 145.115 1.675 145.245 ;
		RECT	1.92 145.115 1.97 145.245 ;
		RECT	5.05 145.115 5.1 145.245 ;
		RECT	1.625 144.655 1.675 144.785 ;
		RECT	1.92 144.655 1.97 144.785 ;
		RECT	5.05 144.655 5.1 144.785 ;
		RECT	3.6 144.195 3.65 144.325 ;
		RECT	1.625 142.235 1.675 142.365 ;
		RECT	1.92 142.235 1.97 142.365 ;
		RECT	5.05 142.235 5.1 142.365 ;
		RECT	1.625 141.775 1.675 141.905 ;
		RECT	1.92 141.775 1.97 141.905 ;
		RECT	5.05 141.775 5.1 141.905 ;
		RECT	3.6 141.315 3.65 141.445 ;
		RECT	1.625 139.355 1.675 139.485 ;
		RECT	1.92 139.355 1.97 139.485 ;
		RECT	5.05 139.355 5.1 139.485 ;
		RECT	1.625 138.895 1.675 139.025 ;
		RECT	1.92 138.895 1.97 139.025 ;
		RECT	5.05 138.895 5.1 139.025 ;
		RECT	3.6 138.435 3.65 138.565 ;
		RECT	1.625 136.475 1.675 136.605 ;
		RECT	1.92 136.475 1.97 136.605 ;
		RECT	5.05 136.475 5.1 136.605 ;
		RECT	1.625 136.015 1.675 136.145 ;
		RECT	1.92 136.015 1.97 136.145 ;
		RECT	5.05 136.015 5.1 136.145 ;
		RECT	3.6 135.555 3.65 135.685 ;
		RECT	1.625 133.595 1.675 133.725 ;
		RECT	1.92 133.595 1.97 133.725 ;
		RECT	5.05 133.595 5.1 133.725 ;
		RECT	1.625 133.135 1.675 133.265 ;
		RECT	1.92 133.135 1.97 133.265 ;
		RECT	5.05 133.135 5.1 133.265 ;
		RECT	3.6 132.675 3.65 132.805 ;
		RECT	1.625 130.715 1.675 130.845 ;
		RECT	1.92 130.715 1.97 130.845 ;
		RECT	5.05 130.715 5.1 130.845 ;
		RECT	1.625 130.255 1.675 130.385 ;
		RECT	1.92 130.255 1.97 130.385 ;
		RECT	5.05 130.255 5.1 130.385 ;
		RECT	3.6 129.795 3.65 129.925 ;
		RECT	1.625 127.835 1.675 127.965 ;
		RECT	1.92 127.835 1.97 127.965 ;
		RECT	5.05 127.835 5.1 127.965 ;
		RECT	1.625 182.095 1.675 182.225 ;
		RECT	1.92 182.095 1.97 182.225 ;
		RECT	5.05 182.095 5.1 182.225 ;
		RECT	3.6 181.635 3.65 181.765 ;
		RECT	1.625 179.675 1.675 179.805 ;
		RECT	1.92 179.675 1.97 179.805 ;
		RECT	5.05 179.675 5.1 179.805 ;
		RECT	1.625 127.375 1.675 127.505 ;
		RECT	1.92 127.375 1.97 127.505 ;
		RECT	5.05 127.375 5.1 127.505 ;
		RECT	3.6 126.915 3.65 127.045 ;
		RECT	1.625 124.955 1.675 125.085 ;
		RECT	1.92 124.955 1.97 125.085 ;
		RECT	5.05 124.955 5.1 125.085 ;
		RECT	1.625 124.495 1.675 124.625 ;
		RECT	1.92 124.495 1.97 124.625 ;
		RECT	5.05 124.495 5.1 124.625 ;
		RECT	3.6 124.035 3.65 124.165 ;
		RECT	1.625 122.075 1.675 122.205 ;
		RECT	1.92 122.075 1.97 122.205 ;
		RECT	5.05 122.075 5.1 122.205 ;
		RECT	1.625 121.615 1.675 121.745 ;
		RECT	1.92 121.615 1.97 121.745 ;
		RECT	5.05 121.615 5.1 121.745 ;
		RECT	3.6 121.155 3.65 121.285 ;
		RECT	1.625 119.195 1.675 119.325 ;
		RECT	1.92 119.195 1.97 119.325 ;
		RECT	5.05 119.195 5.1 119.325 ;
		RECT	1.625 118.735 1.675 118.865 ;
		RECT	1.92 118.735 1.97 118.865 ;
		RECT	5.05 118.735 5.1 118.865 ;
		RECT	3.6 118.275 3.65 118.405 ;
		RECT	1.625 116.315 1.675 116.445 ;
		RECT	1.92 116.315 1.97 116.445 ;
		RECT	5.05 116.315 5.1 116.445 ;
		RECT	1.625 115.855 1.675 115.985 ;
		RECT	1.92 115.855 1.97 115.985 ;
		RECT	5.05 115.855 5.1 115.985 ;
		RECT	3.6 115.395 3.65 115.525 ;
		RECT	1.625 113.435 1.675 113.565 ;
		RECT	1.92 113.435 1.97 113.565 ;
		RECT	5.05 113.435 5.1 113.565 ;
		RECT	1.625 112.975 1.675 113.105 ;
		RECT	1.92 112.975 1.97 113.105 ;
		RECT	5.05 112.975 5.1 113.105 ;
		RECT	3.6 112.515 3.65 112.645 ;
		RECT	1.625 110.555 1.675 110.685 ;
		RECT	1.92 110.555 1.97 110.685 ;
		RECT	5.05 110.555 5.1 110.685 ;
		RECT	1.625 110.095 1.675 110.225 ;
		RECT	1.92 110.095 1.97 110.225 ;
		RECT	5.05 110.095 5.1 110.225 ;
		RECT	3.6 109.635 3.65 109.765 ;
		RECT	1.625 107.675 1.675 107.805 ;
		RECT	1.92 107.675 1.97 107.805 ;
		RECT	5.05 107.675 5.1 107.805 ;
		RECT	1.625 107.215 1.675 107.345 ;
		RECT	1.92 107.215 1.97 107.345 ;
		RECT	5.05 107.215 5.1 107.345 ;
		RECT	3.6 106.755 3.65 106.885 ;
		RECT	1.625 104.795 1.675 104.925 ;
		RECT	1.92 104.795 1.97 104.925 ;
		RECT	5.05 104.795 5.1 104.925 ;
		RECT	1.625 104.335 1.675 104.465 ;
		RECT	1.92 104.335 1.97 104.465 ;
		RECT	5.05 104.335 5.1 104.465 ;
		RECT	3.6 103.875 3.65 104.005 ;
		RECT	1.625 101.915 1.675 102.045 ;
		RECT	1.92 101.915 1.97 102.045 ;
		RECT	5.05 101.915 5.1 102.045 ;
		RECT	1.625 101.455 1.675 101.585 ;
		RECT	1.92 101.455 1.97 101.585 ;
		RECT	5.05 101.455 5.1 101.585 ;
		RECT	3.6 100.995 3.65 101.125 ;
		RECT	1.625 99.035 1.675 99.165 ;
		RECT	1.92 99.035 1.97 99.165 ;
		RECT	5.05 99.035 5.1 99.165 ;
		RECT	1.625 179.215 1.675 179.345 ;
		RECT	1.92 179.215 1.97 179.345 ;
		RECT	5.05 179.215 5.1 179.345 ;
		RECT	3.6 178.755 3.65 178.885 ;
		RECT	1.625 176.795 1.675 176.925 ;
		RECT	1.92 176.795 1.97 176.925 ;
		RECT	5.05 176.795 5.1 176.925 ;
		RECT	1.625 98.575 1.675 98.705 ;
		RECT	1.92 98.575 1.97 98.705 ;
		RECT	5.05 98.575 5.1 98.705 ;
		RECT	3.6 98.115 3.65 98.245 ;
		RECT	1.625 96.155 1.675 96.285 ;
		RECT	1.92 96.155 1.97 96.285 ;
		RECT	5.05 96.155 5.1 96.285 ;
		RECT	1.625 95.695 1.675 95.825 ;
		RECT	1.92 95.695 1.97 95.825 ;
		RECT	5.05 95.695 5.1 95.825 ;
		RECT	3.6 95.235 3.65 95.365 ;
		RECT	1.625 93.275 1.675 93.405 ;
		RECT	1.92 93.275 1.97 93.405 ;
		RECT	5.05 93.275 5.1 93.405 ;
		RECT	1.625 92.815 1.675 92.945 ;
		RECT	1.92 92.815 1.97 92.945 ;
		RECT	5.05 92.815 5.1 92.945 ;
		RECT	3.6 92.355 3.65 92.485 ;
		RECT	1.625 90.395 1.675 90.525 ;
		RECT	1.92 90.395 1.97 90.525 ;
		RECT	5.05 90.395 5.1 90.525 ;
		RECT	1.625 89.935 1.675 90.065 ;
		RECT	1.92 89.935 1.97 90.065 ;
		RECT	5.05 89.935 5.1 90.065 ;
		RECT	3.6 89.475 3.65 89.605 ;
		RECT	1.625 87.515 1.675 87.645 ;
		RECT	1.92 87.515 1.97 87.645 ;
		RECT	5.05 87.515 5.1 87.645 ;
		RECT	1.625 87.055 1.675 87.185 ;
		RECT	1.92 87.055 1.97 87.185 ;
		RECT	5.05 87.055 5.1 87.185 ;
		RECT	3.6 86.595 3.65 86.725 ;
		RECT	1.625 84.635 1.675 84.765 ;
		RECT	1.92 84.635 1.97 84.765 ;
		RECT	5.05 84.635 5.1 84.765 ;
		RECT	1.625 84.175 1.675 84.305 ;
		RECT	1.92 84.175 1.97 84.305 ;
		RECT	5.05 84.175 5.1 84.305 ;
		RECT	3.6 83.715 3.65 83.845 ;
		RECT	1.625 81.755 1.675 81.885 ;
		RECT	1.92 81.755 1.97 81.885 ;
		RECT	5.05 81.755 5.1 81.885 ;
		RECT	1.625 81.295 1.675 81.425 ;
		RECT	1.92 81.295 1.97 81.425 ;
		RECT	5.05 81.295 5.1 81.425 ;
		RECT	3.6 80.835 3.65 80.965 ;
		RECT	1.625 78.875 1.675 79.005 ;
		RECT	1.92 78.875 1.97 79.005 ;
		RECT	5.05 78.875 5.1 79.005 ;
		RECT	1.625 78.415 1.675 78.545 ;
		RECT	1.92 78.415 1.97 78.545 ;
		RECT	5.05 78.415 5.1 78.545 ;
		RECT	3.6 77.955 3.65 78.085 ;
		RECT	1.625 75.995 1.675 76.125 ;
		RECT	1.92 75.995 1.97 76.125 ;
		RECT	5.05 75.995 5.1 76.125 ;
		RECT	1.625 75.535 1.675 75.665 ;
		RECT	1.92 75.535 1.97 75.665 ;
		RECT	5.05 75.535 5.1 75.665 ;
		RECT	3.6 75.075 3.65 75.205 ;
		RECT	1.625 73.115 1.675 73.245 ;
		RECT	1.92 73.115 1.97 73.245 ;
		RECT	5.05 73.115 5.1 73.245 ;
		RECT	1.625 72.655 1.675 72.785 ;
		RECT	1.92 72.655 1.97 72.785 ;
		RECT	5.05 72.655 5.1 72.785 ;
		RECT	3.6 72.195 3.65 72.325 ;
		RECT	1.625 70.235 1.675 70.365 ;
		RECT	1.92 70.235 1.97 70.365 ;
		RECT	5.05 70.235 5.1 70.365 ;
		RECT	1.625 176.335 1.675 176.465 ;
		RECT	1.92 176.335 1.97 176.465 ;
		RECT	5.05 176.335 5.1 176.465 ;
		RECT	3.6 175.875 3.65 176.005 ;
		RECT	1.625 173.915 1.675 174.045 ;
		RECT	1.92 173.915 1.97 174.045 ;
		RECT	5.05 173.915 5.1 174.045 ;
		RECT	1.625 69.775 1.675 69.905 ;
		RECT	1.92 69.775 1.97 69.905 ;
		RECT	5.05 69.775 5.1 69.905 ;
		RECT	3.6 69.315 3.65 69.445 ;
		RECT	1.625 67.355 1.675 67.485 ;
		RECT	1.92 67.355 1.97 67.485 ;
		RECT	5.05 67.355 5.1 67.485 ;
		RECT	1.625 66.895 1.675 67.025 ;
		RECT	1.92 66.895 1.97 67.025 ;
		RECT	5.05 66.895 5.1 67.025 ;
		RECT	3.6 66.435 3.65 66.565 ;
		RECT	1.625 64.475 1.675 64.605 ;
		RECT	1.92 64.475 1.97 64.605 ;
		RECT	5.05 64.475 5.1 64.605 ;
		RECT	1.625 64.015 1.675 64.145 ;
		RECT	1.92 64.015 1.97 64.145 ;
		RECT	5.05 64.015 5.1 64.145 ;
		RECT	3.6 63.555 3.65 63.685 ;
		RECT	1.625 61.595 1.675 61.725 ;
		RECT	1.92 61.595 1.97 61.725 ;
		RECT	5.05 61.595 5.1 61.725 ;
		RECT	1.625 61.135 1.675 61.265 ;
		RECT	1.92 61.135 1.97 61.265 ;
		RECT	5.05 61.135 5.1 61.265 ;
		RECT	3.6 60.675 3.65 60.805 ;
		RECT	1.625 58.715 1.675 58.845 ;
		RECT	1.92 58.715 1.97 58.845 ;
		RECT	5.05 58.715 5.1 58.845 ;
		RECT	1.625 58.255 1.675 58.385 ;
		RECT	1.92 58.255 1.97 58.385 ;
		RECT	5.05 58.255 5.1 58.385 ;
		RECT	3.6 57.795 3.65 57.925 ;
		RECT	1.625 55.835 1.675 55.965 ;
		RECT	1.92 55.835 1.97 55.965 ;
		RECT	5.05 55.835 5.1 55.965 ;
		RECT	1.625 55.375 1.675 55.505 ;
		RECT	1.92 55.375 1.97 55.505 ;
		RECT	5.05 55.375 5.1 55.505 ;
		RECT	3.6 54.915 3.65 55.045 ;
		RECT	1.625 52.955 1.675 53.085 ;
		RECT	1.92 52.955 1.97 53.085 ;
		RECT	5.05 52.955 5.1 53.085 ;
		RECT	1.625 52.495 1.675 52.625 ;
		RECT	1.92 52.495 1.97 52.625 ;
		RECT	5.05 52.495 5.1 52.625 ;
		RECT	3.6 52.035 3.65 52.165 ;
		RECT	1.625 50.075 1.675 50.205 ;
		RECT	1.92 50.075 1.97 50.205 ;
		RECT	5.05 50.075 5.1 50.205 ;
		RECT	1.625 49.615 1.675 49.745 ;
		RECT	1.92 49.615 1.97 49.745 ;
		RECT	5.05 49.615 5.1 49.745 ;
		RECT	3.6 49.155 3.65 49.285 ;
		RECT	1.625 47.195 1.675 47.325 ;
		RECT	1.92 47.195 1.97 47.325 ;
		RECT	5.05 47.195 5.1 47.325 ;
		RECT	1.625 46.735 1.675 46.865 ;
		RECT	1.92 46.735 1.97 46.865 ;
		RECT	5.05 46.735 5.1 46.865 ;
		RECT	3.6 46.275 3.65 46.405 ;
		RECT	1.625 44.315 1.675 44.445 ;
		RECT	1.92 44.315 1.97 44.445 ;
		RECT	5.05 44.315 5.1 44.445 ;
		RECT	1.625 43.855 1.675 43.985 ;
		RECT	1.92 43.855 1.97 43.985 ;
		RECT	5.05 43.855 5.1 43.985 ;
		RECT	3.6 43.395 3.65 43.525 ;
		RECT	1.625 41.435 1.675 41.565 ;
		RECT	1.92 41.435 1.97 41.565 ;
		RECT	5.05 41.435 5.1 41.565 ;
		RECT	1.625 173.455 1.675 173.585 ;
		RECT	1.92 173.455 1.97 173.585 ;
		RECT	5.05 173.455 5.1 173.585 ;
		RECT	3.6 172.995 3.65 173.125 ;
		RECT	1.625 171.035 1.675 171.165 ;
		RECT	1.92 171.035 1.97 171.165 ;
		RECT	5.05 171.035 5.1 171.165 ;
		RECT	1.625 40.975 1.675 41.105 ;
		RECT	1.92 40.975 1.97 41.105 ;
		RECT	5.05 40.975 5.1 41.105 ;
		RECT	3.6 40.515 3.65 40.645 ;
		RECT	1.625 38.555 1.675 38.685 ;
		RECT	1.92 38.555 1.97 38.685 ;
		RECT	5.05 38.555 5.1 38.685 ;
		RECT	1.625 38.095 1.675 38.225 ;
		RECT	1.92 38.095 1.97 38.225 ;
		RECT	5.05 38.095 5.1 38.225 ;
		RECT	3.6 37.635 3.65 37.765 ;
		RECT	1.625 35.675 1.675 35.805 ;
		RECT	1.92 35.675 1.97 35.805 ;
		RECT	5.05 35.675 5.1 35.805 ;
		RECT	1.625 35.215 1.675 35.345 ;
		RECT	1.92 35.215 1.97 35.345 ;
		RECT	5.05 35.215 5.1 35.345 ;
		RECT	3.6 34.755 3.65 34.885 ;
		RECT	1.625 32.795 1.675 32.925 ;
		RECT	1.92 32.795 1.97 32.925 ;
		RECT	5.05 32.795 5.1 32.925 ;
		RECT	1.625 32.335 1.675 32.465 ;
		RECT	1.92 32.335 1.97 32.465 ;
		RECT	5.05 32.335 5.1 32.465 ;
		RECT	3.6 31.875 3.65 32.005 ;
		RECT	1.625 29.915 1.675 30.045 ;
		RECT	1.92 29.915 1.97 30.045 ;
		RECT	5.05 29.915 5.1 30.045 ;
		RECT	1.625 29.455 1.675 29.585 ;
		RECT	1.92 29.455 1.97 29.585 ;
		RECT	5.05 29.455 5.1 29.585 ;
		RECT	3.6 28.995 3.65 29.125 ;
		RECT	1.625 27.035 1.675 27.165 ;
		RECT	1.92 27.035 1.97 27.165 ;
		RECT	5.05 27.035 5.1 27.165 ;
		RECT	1.625 26.575 1.675 26.705 ;
		RECT	1.92 26.575 1.97 26.705 ;
		RECT	5.05 26.575 5.1 26.705 ;
		RECT	3.6 26.115 3.65 26.245 ;
		RECT	1.625 24.155 1.675 24.285 ;
		RECT	1.92 24.155 1.97 24.285 ;
		RECT	5.05 24.155 5.1 24.285 ;
		RECT	1.625 23.695 1.675 23.825 ;
		RECT	1.92 23.695 1.97 23.825 ;
		RECT	5.05 23.695 5.1 23.825 ;
		RECT	3.6 23.235 3.65 23.365 ;
		RECT	1.625 21.275 1.675 21.405 ;
		RECT	1.92 21.275 1.97 21.405 ;
		RECT	5.05 21.275 5.1 21.405 ;
		RECT	1.625 20.815 1.675 20.945 ;
		RECT	1.92 20.815 1.97 20.945 ;
		RECT	5.05 20.815 5.1 20.945 ;
		RECT	3.6 20.355 3.65 20.485 ;
		RECT	1.625 18.395 1.675 18.525 ;
		RECT	1.92 18.395 1.97 18.525 ;
		RECT	5.05 18.395 5.1 18.525 ;
		RECT	1.625 17.935 1.675 18.065 ;
		RECT	1.92 17.935 1.97 18.065 ;
		RECT	5.05 17.935 5.1 18.065 ;
		RECT	3.6 17.475 3.65 17.605 ;
		RECT	1.625 15.515 1.675 15.645 ;
		RECT	1.92 15.515 1.97 15.645 ;
		RECT	5.05 15.515 5.1 15.645 ;
		RECT	1.625 15.055 1.675 15.185 ;
		RECT	1.92 15.055 1.97 15.185 ;
		RECT	5.05 15.055 5.1 15.185 ;
		RECT	3.6 14.595 3.65 14.725 ;
		RECT	1.625 12.635 1.675 12.765 ;
		RECT	1.92 12.635 1.97 12.765 ;
		RECT	5.05 12.635 5.1 12.765 ;
		RECT	1.625 170.575 1.675 170.705 ;
		RECT	1.92 170.575 1.97 170.705 ;
		RECT	5.05 170.575 5.1 170.705 ;
		RECT	3.6 170.115 3.65 170.245 ;
		RECT	1.625 168.155 1.675 168.285 ;
		RECT	1.92 168.155 1.97 168.285 ;
		RECT	5.05 168.155 5.1 168.285 ;
		RECT	1.625 12.175 1.675 12.305 ;
		RECT	1.92 12.175 1.97 12.305 ;
		RECT	5.05 12.175 5.1 12.305 ;
		RECT	3.6 11.715 3.65 11.845 ;
		RECT	1.625 9.755 1.675 9.885 ;
		RECT	1.92 9.755 1.97 9.885 ;
		RECT	5.05 9.755 5.1 9.885 ;
		RECT	1.625 9.295 1.675 9.425 ;
		RECT	1.92 9.295 1.97 9.425 ;
		RECT	5.05 9.295 5.1 9.425 ;
		RECT	3.6 8.835 3.65 8.965 ;
		RECT	1.625 6.875 1.675 7.005 ;
		RECT	1.92 6.875 1.97 7.005 ;
		RECT	5.05 6.875 5.1 7.005 ;
		RECT	1.625 6.415 1.675 6.545 ;
		RECT	1.92 6.415 1.97 6.545 ;
		RECT	5.05 6.415 5.1 6.545 ;
		RECT	3.6 5.955 3.65 6.085 ;
		RECT	1.625 3.995 1.675 4.125 ;
		RECT	1.92 3.995 1.97 4.125 ;
		RECT	5.05 3.995 5.1 4.125 ;
		RECT	1.625 3.535 1.675 3.665 ;
		RECT	1.92 3.535 1.97 3.665 ;
		RECT	5.05 3.535 5.1 3.665 ;
		RECT	3.6 3.075 3.65 3.205 ;
		RECT	1.625 1.115 1.675 1.245 ;
		RECT	1.92 1.115 1.97 1.245 ;
		RECT	5.05 1.115 5.1 1.245 ;
		RECT	1.625 167.695 1.675 167.825 ;
		RECT	1.92 167.695 1.97 167.825 ;
		RECT	5.05 167.695 5.1 167.825 ;
		RECT	3.6 167.235 3.65 167.365 ;
		RECT	1.625 165.275 1.675 165.405 ;
		RECT	1.92 165.275 1.97 165.405 ;
		RECT	5.05 165.275 5.1 165.405 ;
		RECT	1.625 164.815 1.675 164.945 ;
		RECT	1.92 164.815 1.97 164.945 ;
		RECT	5.05 164.815 5.1 164.945 ;
		RECT	3.6 164.355 3.65 164.485 ;
		RECT	1.625 162.395 1.675 162.525 ;
		RECT	1.92 162.395 1.97 162.525 ;
		RECT	5.05 162.395 5.1 162.525 ;
		RECT	1.625 161.935 1.675 162.065 ;
		RECT	1.92 161.935 1.97 162.065 ;
		RECT	5.05 161.935 5.1 162.065 ;
		RECT	3.6 161.475 3.65 161.605 ;
		RECT	1.625 159.515 1.675 159.645 ;
		RECT	1.92 159.515 1.97 159.645 ;
		RECT	5.05 159.515 5.1 159.645 ;
		RECT	1.625 159.055 1.675 159.185 ;
		RECT	1.92 159.055 1.97 159.185 ;
		RECT	5.05 159.055 5.1 159.185 ;
		RECT	3.6 158.595 3.65 158.725 ;
		RECT	1.625 156.635 1.675 156.765 ;
		RECT	1.92 156.635 1.97 156.765 ;
		RECT	5.05 156.635 5.1 156.765 ;
		RECT	3.6 182.095 3.65 182.225 ;
		RECT	1.625 181.635 1.675 181.765 ;
		RECT	1.88 181.675 2.01 181.725 ;
		RECT	5.01 181.675 5.14 181.725 ;
		RECT	3.6 179.675 3.65 179.805 ;
		RECT	1.44 179.445 1.49 179.575 ;
		RECT	2.11 179.445 2.16 179.575 ;
		RECT	3.09 179.445 3.14 179.575 ;
		RECT	4.38 179.445 4.43 179.575 ;
		RECT	6.215 179.445 6.265 179.575 ;
		RECT	3.6 156.175 3.65 156.305 ;
		RECT	1.625 155.715 1.675 155.845 ;
		RECT	1.88 155.755 2.01 155.805 ;
		RECT	5.01 155.755 5.14 155.805 ;
		RECT	3.6 153.755 3.65 153.885 ;
		RECT	1.44 153.525 1.49 153.655 ;
		RECT	2.11 153.525 2.16 153.655 ;
		RECT	3.09 153.525 3.14 153.655 ;
		RECT	4.38 153.525 4.43 153.655 ;
		RECT	6.215 153.525 6.265 153.655 ;
		RECT	3.6 153.295 3.65 153.425 ;
		RECT	1.625 152.835 1.675 152.965 ;
		RECT	1.88 152.875 2.01 152.925 ;
		RECT	5.01 152.875 5.14 152.925 ;
		RECT	3.6 150.875 3.65 151.005 ;
		RECT	1.44 150.645 1.49 150.775 ;
		RECT	2.11 150.645 2.16 150.775 ;
		RECT	3.09 150.645 3.14 150.775 ;
		RECT	4.38 150.645 4.43 150.775 ;
		RECT	6.215 150.645 6.265 150.775 ;
		RECT	3.6 150.415 3.65 150.545 ;
		RECT	1.625 149.955 1.675 150.085 ;
		RECT	1.88 149.995 2.01 150.045 ;
		RECT	5.01 149.995 5.14 150.045 ;
		RECT	3.6 147.995 3.65 148.125 ;
		RECT	1.44 147.765 1.49 147.895 ;
		RECT	2.11 147.765 2.16 147.895 ;
		RECT	3.09 147.765 3.14 147.895 ;
		RECT	4.38 147.765 4.43 147.895 ;
		RECT	6.215 147.765 6.265 147.895 ;
		RECT	3.6 147.535 3.65 147.665 ;
		RECT	1.625 147.075 1.675 147.205 ;
		RECT	1.88 147.115 2.01 147.165 ;
		RECT	5.01 147.115 5.14 147.165 ;
		RECT	3.6 145.115 3.65 145.245 ;
		RECT	1.44 144.885 1.49 145.015 ;
		RECT	2.11 144.885 2.16 145.015 ;
		RECT	3.09 144.885 3.14 145.015 ;
		RECT	4.38 144.885 4.43 145.015 ;
		RECT	6.215 144.885 6.265 145.015 ;
		RECT	3.6 144.655 3.65 144.785 ;
		RECT	1.625 144.195 1.675 144.325 ;
		RECT	1.88 144.235 2.01 144.285 ;
		RECT	5.01 144.235 5.14 144.285 ;
		RECT	3.6 142.235 3.65 142.365 ;
		RECT	1.44 142.005 1.49 142.135 ;
		RECT	2.11 142.005 2.16 142.135 ;
		RECT	3.09 142.005 3.14 142.135 ;
		RECT	4.38 142.005 4.43 142.135 ;
		RECT	6.215 142.005 6.265 142.135 ;
		RECT	3.6 141.775 3.65 141.905 ;
		RECT	1.625 141.315 1.675 141.445 ;
		RECT	1.88 141.355 2.01 141.405 ;
		RECT	5.01 141.355 5.14 141.405 ;
		RECT	3.6 139.355 3.65 139.485 ;
		RECT	1.44 139.125 1.49 139.255 ;
		RECT	2.11 139.125 2.16 139.255 ;
		RECT	3.09 139.125 3.14 139.255 ;
		RECT	4.38 139.125 4.43 139.255 ;
		RECT	6.215 139.125 6.265 139.255 ;
		RECT	3.6 138.895 3.65 139.025 ;
		RECT	1.625 138.435 1.675 138.565 ;
		RECT	1.88 138.475 2.01 138.525 ;
		RECT	5.01 138.475 5.14 138.525 ;
		RECT	3.6 136.475 3.65 136.605 ;
		RECT	1.44 136.245 1.49 136.375 ;
		RECT	2.11 136.245 2.16 136.375 ;
		RECT	3.09 136.245 3.14 136.375 ;
		RECT	4.38 136.245 4.43 136.375 ;
		RECT	6.215 136.245 6.265 136.375 ;
		RECT	3.6 136.015 3.65 136.145 ;
		RECT	1.625 135.555 1.675 135.685 ;
		RECT	1.88 135.595 2.01 135.645 ;
		RECT	5.01 135.595 5.14 135.645 ;
		RECT	3.6 133.595 3.65 133.725 ;
		RECT	1.44 133.365 1.49 133.495 ;
		RECT	2.11 133.365 2.16 133.495 ;
		RECT	3.09 133.365 3.14 133.495 ;
		RECT	4.38 133.365 4.43 133.495 ;
		RECT	6.215 133.365 6.265 133.495 ;
		RECT	3.6 133.135 3.65 133.265 ;
		RECT	1.625 132.675 1.675 132.805 ;
		RECT	1.88 132.715 2.01 132.765 ;
		RECT	5.01 132.715 5.14 132.765 ;
		RECT	3.6 130.715 3.65 130.845 ;
		RECT	1.44 130.485 1.49 130.615 ;
		RECT	2.11 130.485 2.16 130.615 ;
		RECT	3.09 130.485 3.14 130.615 ;
		RECT	4.38 130.485 4.43 130.615 ;
		RECT	6.215 130.485 6.265 130.615 ;
		RECT	3.6 130.255 3.65 130.385 ;
		RECT	1.625 129.795 1.675 129.925 ;
		RECT	1.88 129.835 2.01 129.885 ;
		RECT	5.01 129.835 5.14 129.885 ;
		RECT	3.6 127.835 3.65 127.965 ;
		RECT	1.44 127.605 1.49 127.735 ;
		RECT	2.11 127.605 2.16 127.735 ;
		RECT	3.09 127.605 3.14 127.735 ;
		RECT	4.38 127.605 4.43 127.735 ;
		RECT	6.215 127.605 6.265 127.735 ;
		RECT	3.6 179.215 3.65 179.345 ;
		RECT	1.625 178.755 1.675 178.885 ;
		RECT	1.88 178.795 2.01 178.845 ;
		RECT	5.01 178.795 5.14 178.845 ;
		RECT	3.6 176.795 3.65 176.925 ;
		RECT	1.44 176.565 1.49 176.695 ;
		RECT	2.11 176.565 2.16 176.695 ;
		RECT	3.09 176.565 3.14 176.695 ;
		RECT	4.38 176.565 4.43 176.695 ;
		RECT	6.215 176.565 6.265 176.695 ;
		RECT	3.6 127.375 3.65 127.505 ;
		RECT	1.625 126.915 1.675 127.045 ;
		RECT	1.88 126.955 2.01 127.005 ;
		RECT	5.01 126.955 5.14 127.005 ;
		RECT	3.6 124.955 3.65 125.085 ;
		RECT	1.44 124.725 1.49 124.855 ;
		RECT	2.11 124.725 2.16 124.855 ;
		RECT	3.09 124.725 3.14 124.855 ;
		RECT	4.38 124.725 4.43 124.855 ;
		RECT	6.215 124.725 6.265 124.855 ;
		RECT	3.6 124.495 3.65 124.625 ;
		RECT	1.625 124.035 1.675 124.165 ;
		RECT	1.88 124.075 2.01 124.125 ;
		RECT	5.01 124.075 5.14 124.125 ;
		RECT	3.6 122.075 3.65 122.205 ;
		RECT	1.44 121.845 1.49 121.975 ;
		RECT	2.11 121.845 2.16 121.975 ;
		RECT	3.09 121.845 3.14 121.975 ;
		RECT	4.38 121.845 4.43 121.975 ;
		RECT	6.215 121.845 6.265 121.975 ;
		RECT	3.6 121.615 3.65 121.745 ;
		RECT	1.625 121.155 1.675 121.285 ;
		RECT	1.88 121.195 2.01 121.245 ;
		RECT	5.01 121.195 5.14 121.245 ;
		RECT	3.6 119.195 3.65 119.325 ;
		RECT	1.44 118.965 1.49 119.095 ;
		RECT	2.11 118.965 2.16 119.095 ;
		RECT	3.09 118.965 3.14 119.095 ;
		RECT	4.38 118.965 4.43 119.095 ;
		RECT	6.215 118.965 6.265 119.095 ;
		RECT	3.6 118.735 3.65 118.865 ;
		RECT	1.625 118.275 1.675 118.405 ;
		RECT	1.88 118.315 2.01 118.365 ;
		RECT	5.01 118.315 5.14 118.365 ;
		RECT	3.6 116.315 3.65 116.445 ;
		RECT	1.44 116.085 1.49 116.215 ;
		RECT	2.11 116.085 2.16 116.215 ;
		RECT	3.09 116.085 3.14 116.215 ;
		RECT	4.38 116.085 4.43 116.215 ;
		RECT	6.215 116.085 6.265 116.215 ;
		RECT	3.6 115.855 3.65 115.985 ;
		RECT	1.625 115.395 1.675 115.525 ;
		RECT	1.88 115.435 2.01 115.485 ;
		RECT	5.01 115.435 5.14 115.485 ;
		RECT	3.6 113.435 3.65 113.565 ;
		RECT	1.44 113.205 1.49 113.335 ;
		RECT	2.11 113.205 2.16 113.335 ;
		RECT	3.09 113.205 3.14 113.335 ;
		RECT	4.38 113.205 4.43 113.335 ;
		RECT	6.215 113.205 6.265 113.335 ;
		RECT	3.6 112.975 3.65 113.105 ;
		RECT	1.625 112.515 1.675 112.645 ;
		RECT	1.88 112.555 2.01 112.605 ;
		RECT	5.01 112.555 5.14 112.605 ;
		RECT	3.6 110.555 3.65 110.685 ;
		RECT	1.44 110.325 1.49 110.455 ;
		RECT	2.11 110.325 2.16 110.455 ;
		RECT	3.09 110.325 3.14 110.455 ;
		RECT	4.38 110.325 4.43 110.455 ;
		RECT	6.215 110.325 6.265 110.455 ;
		RECT	3.6 110.095 3.65 110.225 ;
		RECT	1.625 109.635 1.675 109.765 ;
		RECT	1.88 109.675 2.01 109.725 ;
		RECT	5.01 109.675 5.14 109.725 ;
		RECT	3.6 107.675 3.65 107.805 ;
		RECT	1.44 107.445 1.49 107.575 ;
		RECT	2.11 107.445 2.16 107.575 ;
		RECT	3.09 107.445 3.14 107.575 ;
		RECT	4.38 107.445 4.43 107.575 ;
		RECT	6.215 107.445 6.265 107.575 ;
		RECT	3.6 107.215 3.65 107.345 ;
		RECT	1.625 106.755 1.675 106.885 ;
		RECT	1.88 106.795 2.01 106.845 ;
		RECT	5.01 106.795 5.14 106.845 ;
		RECT	3.6 104.795 3.65 104.925 ;
		RECT	1.44 104.565 1.49 104.695 ;
		RECT	2.11 104.565 2.16 104.695 ;
		RECT	3.09 104.565 3.14 104.695 ;
		RECT	4.38 104.565 4.43 104.695 ;
		RECT	6.215 104.565 6.265 104.695 ;
		RECT	3.6 104.335 3.65 104.465 ;
		RECT	1.625 103.875 1.675 104.005 ;
		RECT	1.88 103.915 2.01 103.965 ;
		RECT	5.01 103.915 5.14 103.965 ;
		RECT	3.6 101.915 3.65 102.045 ;
		RECT	1.44 101.685 1.49 101.815 ;
		RECT	2.11 101.685 2.16 101.815 ;
		RECT	3.09 101.685 3.14 101.815 ;
		RECT	4.38 101.685 4.43 101.815 ;
		RECT	6.215 101.685 6.265 101.815 ;
		RECT	3.6 101.455 3.65 101.585 ;
		RECT	1.625 100.995 1.675 101.125 ;
		RECT	1.88 101.035 2.01 101.085 ;
		RECT	5.01 101.035 5.14 101.085 ;
		RECT	3.6 99.035 3.65 99.165 ;
		RECT	1.44 98.805 1.49 98.935 ;
		RECT	2.11 98.805 2.16 98.935 ;
		RECT	3.09 98.805 3.14 98.935 ;
		RECT	4.38 98.805 4.43 98.935 ;
		RECT	6.215 98.805 6.265 98.935 ;
		RECT	3.6 176.335 3.65 176.465 ;
		RECT	1.625 175.875 1.675 176.005 ;
		RECT	1.88 175.915 2.01 175.965 ;
		RECT	5.01 175.915 5.14 175.965 ;
		RECT	3.6 173.915 3.65 174.045 ;
		RECT	1.44 173.685 1.49 173.815 ;
		RECT	2.11 173.685 2.16 173.815 ;
		RECT	3.09 173.685 3.14 173.815 ;
		RECT	4.38 173.685 4.43 173.815 ;
		RECT	6.215 173.685 6.265 173.815 ;
		RECT	3.6 98.575 3.65 98.705 ;
		RECT	1.625 98.115 1.675 98.245 ;
		RECT	1.88 98.155 2.01 98.205 ;
		RECT	5.01 98.155 5.14 98.205 ;
		RECT	3.6 96.155 3.65 96.285 ;
		RECT	1.44 95.925 1.49 96.055 ;
		RECT	2.11 95.925 2.16 96.055 ;
		RECT	3.09 95.925 3.14 96.055 ;
		RECT	4.38 95.925 4.43 96.055 ;
		RECT	6.215 95.925 6.265 96.055 ;
		RECT	3.6 95.695 3.65 95.825 ;
		RECT	1.625 95.235 1.675 95.365 ;
		RECT	1.88 95.275 2.01 95.325 ;
		RECT	5.01 95.275 5.14 95.325 ;
		RECT	3.6 93.275 3.65 93.405 ;
		RECT	1.44 93.045 1.49 93.175 ;
		RECT	2.11 93.045 2.16 93.175 ;
		RECT	3.09 93.045 3.14 93.175 ;
		RECT	4.38 93.045 4.43 93.175 ;
		RECT	6.215 93.045 6.265 93.175 ;
		RECT	3.6 92.815 3.65 92.945 ;
		RECT	1.625 92.355 1.675 92.485 ;
		RECT	1.88 92.395 2.01 92.445 ;
		RECT	5.01 92.395 5.14 92.445 ;
		RECT	3.6 90.395 3.65 90.525 ;
		RECT	1.44 90.165 1.49 90.295 ;
		RECT	2.11 90.165 2.16 90.295 ;
		RECT	3.09 90.165 3.14 90.295 ;
		RECT	4.38 90.165 4.43 90.295 ;
		RECT	6.215 90.165 6.265 90.295 ;
		RECT	3.6 89.935 3.65 90.065 ;
		RECT	1.625 89.475 1.675 89.605 ;
		RECT	1.88 89.515 2.01 89.565 ;
		RECT	5.01 89.515 5.14 89.565 ;
		RECT	3.6 87.515 3.65 87.645 ;
		RECT	1.44 87.285 1.49 87.415 ;
		RECT	2.11 87.285 2.16 87.415 ;
		RECT	3.09 87.285 3.14 87.415 ;
		RECT	4.38 87.285 4.43 87.415 ;
		RECT	6.215 87.285 6.265 87.415 ;
		RECT	3.6 87.055 3.65 87.185 ;
		RECT	1.625 86.595 1.675 86.725 ;
		RECT	1.88 86.635 2.01 86.685 ;
		RECT	5.01 86.635 5.14 86.685 ;
		RECT	3.6 84.635 3.65 84.765 ;
		RECT	1.44 84.405 1.49 84.535 ;
		RECT	2.11 84.405 2.16 84.535 ;
		RECT	3.09 84.405 3.14 84.535 ;
		RECT	4.38 84.405 4.43 84.535 ;
		RECT	6.215 84.405 6.265 84.535 ;
		RECT	3.6 84.175 3.65 84.305 ;
		RECT	1.625 83.715 1.675 83.845 ;
		RECT	1.88 83.755 2.01 83.805 ;
		RECT	5.01 83.755 5.14 83.805 ;
		RECT	3.6 81.755 3.65 81.885 ;
		RECT	1.44 81.525 1.49 81.655 ;
		RECT	2.11 81.525 2.16 81.655 ;
		RECT	3.09 81.525 3.14 81.655 ;
		RECT	4.38 81.525 4.43 81.655 ;
		RECT	6.215 81.525 6.265 81.655 ;
		RECT	3.6 81.295 3.65 81.425 ;
		RECT	1.625 80.835 1.675 80.965 ;
		RECT	1.88 80.875 2.01 80.925 ;
		RECT	5.01 80.875 5.14 80.925 ;
		RECT	3.6 78.875 3.65 79.005 ;
		RECT	1.44 78.645 1.49 78.775 ;
		RECT	2.11 78.645 2.16 78.775 ;
		RECT	3.09 78.645 3.14 78.775 ;
		RECT	4.38 78.645 4.43 78.775 ;
		RECT	6.215 78.645 6.265 78.775 ;
		RECT	3.6 78.415 3.65 78.545 ;
		RECT	1.625 77.955 1.675 78.085 ;
		RECT	1.88 77.995 2.01 78.045 ;
		RECT	5.01 77.995 5.14 78.045 ;
		RECT	3.6 75.995 3.65 76.125 ;
		RECT	1.44 75.765 1.49 75.895 ;
		RECT	2.11 75.765 2.16 75.895 ;
		RECT	3.09 75.765 3.14 75.895 ;
		RECT	4.38 75.765 4.43 75.895 ;
		RECT	6.215 75.765 6.265 75.895 ;
		RECT	3.6 75.535 3.65 75.665 ;
		RECT	1.625 75.075 1.675 75.205 ;
		RECT	1.88 75.115 2.01 75.165 ;
		RECT	5.01 75.115 5.14 75.165 ;
		RECT	3.6 73.115 3.65 73.245 ;
		RECT	1.44 72.885 1.49 73.015 ;
		RECT	2.11 72.885 2.16 73.015 ;
		RECT	3.09 72.885 3.14 73.015 ;
		RECT	4.38 72.885 4.43 73.015 ;
		RECT	6.215 72.885 6.265 73.015 ;
		RECT	3.6 72.655 3.65 72.785 ;
		RECT	1.625 72.195 1.675 72.325 ;
		RECT	1.88 72.235 2.01 72.285 ;
		RECT	5.01 72.235 5.14 72.285 ;
		RECT	3.6 70.235 3.65 70.365 ;
		RECT	1.44 70.005 1.49 70.135 ;
		RECT	2.11 70.005 2.16 70.135 ;
		RECT	3.09 70.005 3.14 70.135 ;
		RECT	4.38 70.005 4.43 70.135 ;
		RECT	6.215 70.005 6.265 70.135 ;
		RECT	3.6 173.455 3.65 173.585 ;
		RECT	1.625 172.995 1.675 173.125 ;
		RECT	1.88 173.035 2.01 173.085 ;
		RECT	5.01 173.035 5.14 173.085 ;
		RECT	3.6 171.035 3.65 171.165 ;
		RECT	1.44 170.805 1.49 170.935 ;
		RECT	2.11 170.805 2.16 170.935 ;
		RECT	3.09 170.805 3.14 170.935 ;
		RECT	4.38 170.805 4.43 170.935 ;
		RECT	6.215 170.805 6.265 170.935 ;
		RECT	3.6 69.775 3.65 69.905 ;
		RECT	1.625 69.315 1.675 69.445 ;
		RECT	1.88 69.355 2.01 69.405 ;
		RECT	5.01 69.355 5.14 69.405 ;
		RECT	3.6 67.355 3.65 67.485 ;
		RECT	1.44 67.125 1.49 67.255 ;
		RECT	2.11 67.125 2.16 67.255 ;
		RECT	3.09 67.125 3.14 67.255 ;
		RECT	4.38 67.125 4.43 67.255 ;
		RECT	6.215 67.125 6.265 67.255 ;
		RECT	3.6 66.895 3.65 67.025 ;
		RECT	1.625 66.435 1.675 66.565 ;
		RECT	1.88 66.475 2.01 66.525 ;
		RECT	5.01 66.475 5.14 66.525 ;
		RECT	3.6 64.475 3.65 64.605 ;
		RECT	1.44 64.245 1.49 64.375 ;
		RECT	2.11 64.245 2.16 64.375 ;
		RECT	3.09 64.245 3.14 64.375 ;
		RECT	4.38 64.245 4.43 64.375 ;
		RECT	6.215 64.245 6.265 64.375 ;
		RECT	3.6 64.015 3.65 64.145 ;
		RECT	1.625 63.555 1.675 63.685 ;
		RECT	1.88 63.595 2.01 63.645 ;
		RECT	5.01 63.595 5.14 63.645 ;
		RECT	3.6 61.595 3.65 61.725 ;
		RECT	1.44 61.365 1.49 61.495 ;
		RECT	2.11 61.365 2.16 61.495 ;
		RECT	3.09 61.365 3.14 61.495 ;
		RECT	4.38 61.365 4.43 61.495 ;
		RECT	6.215 61.365 6.265 61.495 ;
		RECT	3.6 61.135 3.65 61.265 ;
		RECT	1.625 60.675 1.675 60.805 ;
		RECT	1.88 60.715 2.01 60.765 ;
		RECT	5.01 60.715 5.14 60.765 ;
		RECT	3.6 58.715 3.65 58.845 ;
		RECT	1.44 58.485 1.49 58.615 ;
		RECT	2.11 58.485 2.16 58.615 ;
		RECT	3.09 58.485 3.14 58.615 ;
		RECT	4.38 58.485 4.43 58.615 ;
		RECT	6.215 58.485 6.265 58.615 ;
		RECT	3.6 58.255 3.65 58.385 ;
		RECT	1.625 57.795 1.675 57.925 ;
		RECT	1.88 57.835 2.01 57.885 ;
		RECT	5.01 57.835 5.14 57.885 ;
		RECT	3.6 55.835 3.65 55.965 ;
		RECT	1.44 55.605 1.49 55.735 ;
		RECT	2.11 55.605 2.16 55.735 ;
		RECT	3.09 55.605 3.14 55.735 ;
		RECT	4.38 55.605 4.43 55.735 ;
		RECT	6.215 55.605 6.265 55.735 ;
		RECT	3.6 55.375 3.65 55.505 ;
		RECT	1.625 54.915 1.675 55.045 ;
		RECT	1.88 54.955 2.01 55.005 ;
		RECT	5.01 54.955 5.14 55.005 ;
		RECT	3.6 52.955 3.65 53.085 ;
		RECT	1.44 52.725 1.49 52.855 ;
		RECT	2.11 52.725 2.16 52.855 ;
		RECT	3.09 52.725 3.14 52.855 ;
		RECT	4.38 52.725 4.43 52.855 ;
		RECT	6.215 52.725 6.265 52.855 ;
		RECT	3.6 52.495 3.65 52.625 ;
		RECT	1.625 52.035 1.675 52.165 ;
		RECT	1.88 52.075 2.01 52.125 ;
		RECT	5.01 52.075 5.14 52.125 ;
		RECT	3.6 50.075 3.65 50.205 ;
		RECT	1.44 49.845 1.49 49.975 ;
		RECT	2.11 49.845 2.16 49.975 ;
		RECT	3.09 49.845 3.14 49.975 ;
		RECT	4.38 49.845 4.43 49.975 ;
		RECT	6.215 49.845 6.265 49.975 ;
		RECT	3.6 49.615 3.65 49.745 ;
		RECT	1.625 49.155 1.675 49.285 ;
		RECT	1.88 49.195 2.01 49.245 ;
		RECT	5.01 49.195 5.14 49.245 ;
		RECT	3.6 47.195 3.65 47.325 ;
		RECT	1.44 46.965 1.49 47.095 ;
		RECT	2.11 46.965 2.16 47.095 ;
		RECT	3.09 46.965 3.14 47.095 ;
		RECT	4.38 46.965 4.43 47.095 ;
		RECT	6.215 46.965 6.265 47.095 ;
		RECT	3.6 46.735 3.65 46.865 ;
		RECT	1.625 46.275 1.675 46.405 ;
		RECT	1.88 46.315 2.01 46.365 ;
		RECT	5.01 46.315 5.14 46.365 ;
		RECT	3.6 44.315 3.65 44.445 ;
		RECT	1.44 44.085 1.49 44.215 ;
		RECT	2.11 44.085 2.16 44.215 ;
		RECT	3.09 44.085 3.14 44.215 ;
		RECT	4.38 44.085 4.43 44.215 ;
		RECT	6.215 44.085 6.265 44.215 ;
		RECT	3.6 43.855 3.65 43.985 ;
		RECT	1.625 43.395 1.675 43.525 ;
		RECT	1.88 43.435 2.01 43.485 ;
		RECT	5.01 43.435 5.14 43.485 ;
		RECT	3.6 41.435 3.65 41.565 ;
		RECT	1.44 41.205 1.49 41.335 ;
		RECT	2.11 41.205 2.16 41.335 ;
		RECT	3.09 41.205 3.14 41.335 ;
		RECT	4.38 41.205 4.43 41.335 ;
		RECT	6.215 41.205 6.265 41.335 ;
		RECT	3.6 170.575 3.65 170.705 ;
		RECT	1.625 170.115 1.675 170.245 ;
		RECT	1.88 170.155 2.01 170.205 ;
		RECT	5.01 170.155 5.14 170.205 ;
		RECT	3.6 168.155 3.65 168.285 ;
		RECT	1.44 167.925 1.49 168.055 ;
		RECT	2.11 167.925 2.16 168.055 ;
		RECT	3.09 167.925 3.14 168.055 ;
		RECT	4.38 167.925 4.43 168.055 ;
		RECT	6.215 167.925 6.265 168.055 ;
		RECT	3.6 40.975 3.65 41.105 ;
		RECT	1.625 40.515 1.675 40.645 ;
		RECT	1.88 40.555 2.01 40.605 ;
		RECT	5.01 40.555 5.14 40.605 ;
		RECT	3.6 38.555 3.65 38.685 ;
		RECT	1.44 38.325 1.49 38.455 ;
		RECT	2.11 38.325 2.16 38.455 ;
		RECT	3.09 38.325 3.14 38.455 ;
		RECT	4.38 38.325 4.43 38.455 ;
		RECT	6.215 38.325 6.265 38.455 ;
		RECT	3.6 38.095 3.65 38.225 ;
		RECT	1.625 37.635 1.675 37.765 ;
		RECT	1.88 37.675 2.01 37.725 ;
		RECT	5.01 37.675 5.14 37.725 ;
		RECT	3.6 35.675 3.65 35.805 ;
		RECT	1.44 35.445 1.49 35.575 ;
		RECT	2.11 35.445 2.16 35.575 ;
		RECT	3.09 35.445 3.14 35.575 ;
		RECT	4.38 35.445 4.43 35.575 ;
		RECT	6.215 35.445 6.265 35.575 ;
		RECT	3.6 35.215 3.65 35.345 ;
		RECT	1.625 34.755 1.675 34.885 ;
		RECT	1.88 34.795 2.01 34.845 ;
		RECT	5.01 34.795 5.14 34.845 ;
		RECT	3.6 32.795 3.65 32.925 ;
		RECT	1.44 32.565 1.49 32.695 ;
		RECT	2.11 32.565 2.16 32.695 ;
		RECT	3.09 32.565 3.14 32.695 ;
		RECT	4.38 32.565 4.43 32.695 ;
		RECT	6.215 32.565 6.265 32.695 ;
		RECT	3.6 32.335 3.65 32.465 ;
		RECT	1.625 31.875 1.675 32.005 ;
		RECT	1.88 31.915 2.01 31.965 ;
		RECT	5.01 31.915 5.14 31.965 ;
		RECT	3.6 29.915 3.65 30.045 ;
		RECT	1.44 29.685 1.49 29.815 ;
		RECT	2.11 29.685 2.16 29.815 ;
		RECT	3.09 29.685 3.14 29.815 ;
		RECT	4.38 29.685 4.43 29.815 ;
		RECT	6.215 29.685 6.265 29.815 ;
		RECT	3.6 29.455 3.65 29.585 ;
		RECT	1.625 28.995 1.675 29.125 ;
		RECT	1.88 29.035 2.01 29.085 ;
		RECT	5.01 29.035 5.14 29.085 ;
		RECT	3.6 27.035 3.65 27.165 ;
		RECT	1.44 26.805 1.49 26.935 ;
		RECT	2.11 26.805 2.16 26.935 ;
		RECT	3.09 26.805 3.14 26.935 ;
		RECT	4.38 26.805 4.43 26.935 ;
		RECT	6.215 26.805 6.265 26.935 ;
		RECT	3.6 26.575 3.65 26.705 ;
		RECT	1.625 26.115 1.675 26.245 ;
		RECT	1.88 26.155 2.01 26.205 ;
		RECT	5.01 26.155 5.14 26.205 ;
		RECT	3.6 24.155 3.65 24.285 ;
		RECT	1.44 23.925 1.49 24.055 ;
		RECT	2.11 23.925 2.16 24.055 ;
		RECT	3.09 23.925 3.14 24.055 ;
		RECT	4.38 23.925 4.43 24.055 ;
		RECT	6.215 23.925 6.265 24.055 ;
		RECT	3.6 23.695 3.65 23.825 ;
		RECT	1.625 23.235 1.675 23.365 ;
		RECT	1.88 23.275 2.01 23.325 ;
		RECT	5.01 23.275 5.14 23.325 ;
		RECT	3.6 21.275 3.65 21.405 ;
		RECT	1.44 21.045 1.49 21.175 ;
		RECT	2.11 21.045 2.16 21.175 ;
		RECT	3.09 21.045 3.14 21.175 ;
		RECT	4.38 21.045 4.43 21.175 ;
		RECT	6.215 21.045 6.265 21.175 ;
		RECT	3.6 20.815 3.65 20.945 ;
		RECT	1.625 20.355 1.675 20.485 ;
		RECT	1.88 20.395 2.01 20.445 ;
		RECT	5.01 20.395 5.14 20.445 ;
		RECT	3.6 18.395 3.65 18.525 ;
		RECT	1.44 18.165 1.49 18.295 ;
		RECT	2.11 18.165 2.16 18.295 ;
		RECT	3.09 18.165 3.14 18.295 ;
		RECT	4.38 18.165 4.43 18.295 ;
		RECT	6.215 18.165 6.265 18.295 ;
		RECT	3.6 17.935 3.65 18.065 ;
		RECT	1.625 17.475 1.675 17.605 ;
		RECT	1.88 17.515 2.01 17.565 ;
		RECT	5.01 17.515 5.14 17.565 ;
		RECT	3.6 15.515 3.65 15.645 ;
		RECT	1.44 15.285 1.49 15.415 ;
		RECT	2.11 15.285 2.16 15.415 ;
		RECT	3.09 15.285 3.14 15.415 ;
		RECT	4.38 15.285 4.43 15.415 ;
		RECT	6.215 15.285 6.265 15.415 ;
		RECT	3.6 15.055 3.65 15.185 ;
		RECT	1.625 14.595 1.675 14.725 ;
		RECT	1.88 14.635 2.01 14.685 ;
		RECT	5.01 14.635 5.14 14.685 ;
		RECT	3.6 12.635 3.65 12.765 ;
		RECT	1.44 12.405 1.49 12.535 ;
		RECT	2.11 12.405 2.16 12.535 ;
		RECT	3.09 12.405 3.14 12.535 ;
		RECT	4.38 12.405 4.43 12.535 ;
		RECT	6.215 12.405 6.265 12.535 ;
		RECT	3.6 167.695 3.65 167.825 ;
		RECT	1.625 167.235 1.675 167.365 ;
		RECT	1.88 167.275 2.01 167.325 ;
		RECT	5.01 167.275 5.14 167.325 ;
		RECT	3.6 165.275 3.65 165.405 ;
		RECT	1.44 165.045 1.49 165.175 ;
		RECT	2.11 165.045 2.16 165.175 ;
		RECT	3.09 165.045 3.14 165.175 ;
		RECT	4.38 165.045 4.43 165.175 ;
		RECT	6.215 165.045 6.265 165.175 ;
		RECT	3.6 12.175 3.65 12.305 ;
		RECT	1.625 11.715 1.675 11.845 ;
		RECT	1.88 11.755 2.01 11.805 ;
		RECT	5.01 11.755 5.14 11.805 ;
		RECT	3.6 9.755 3.65 9.885 ;
		RECT	1.44 9.525 1.49 9.655 ;
		RECT	2.11 9.525 2.16 9.655 ;
		RECT	3.09 9.525 3.14 9.655 ;
		RECT	4.38 9.525 4.43 9.655 ;
		RECT	6.215 9.525 6.265 9.655 ;
		RECT	3.6 9.295 3.65 9.425 ;
		RECT	1.625 8.835 1.675 8.965 ;
		RECT	1.88 8.875 2.01 8.925 ;
		RECT	5.01 8.875 5.14 8.925 ;
		RECT	3.6 6.875 3.65 7.005 ;
		RECT	1.44 6.645 1.49 6.775 ;
		RECT	2.11 6.645 2.16 6.775 ;
		RECT	3.09 6.645 3.14 6.775 ;
		RECT	4.38 6.645 4.43 6.775 ;
		RECT	6.215 6.645 6.265 6.775 ;
		RECT	3.6 6.415 3.65 6.545 ;
		RECT	1.625 5.955 1.675 6.085 ;
		RECT	1.88 5.995 2.01 6.045 ;
		RECT	5.01 5.995 5.14 6.045 ;
		RECT	3.6 3.995 3.65 4.125 ;
		RECT	1.44 3.765 1.49 3.895 ;
		RECT	2.11 3.765 2.16 3.895 ;
		RECT	3.09 3.765 3.14 3.895 ;
		RECT	4.38 3.765 4.43 3.895 ;
		RECT	6.215 3.765 6.265 3.895 ;
		RECT	3.6 164.815 3.65 164.945 ;
		RECT	1.625 164.355 1.675 164.485 ;
		RECT	1.88 164.395 2.01 164.445 ;
		RECT	5.01 164.395 5.14 164.445 ;
		RECT	3.6 162.395 3.65 162.525 ;
		RECT	1.44 162.165 1.49 162.295 ;
		RECT	2.11 162.165 2.16 162.295 ;
		RECT	3.09 162.165 3.14 162.295 ;
		RECT	4.38 162.165 4.43 162.295 ;
		RECT	6.215 162.165 6.265 162.295 ;
		RECT	3.6 161.935 3.65 162.065 ;
		RECT	1.625 161.475 1.675 161.605 ;
		RECT	1.88 161.515 2.01 161.565 ;
		RECT	5.01 161.515 5.14 161.565 ;
		RECT	3.6 159.515 3.65 159.645 ;
		RECT	1.44 159.285 1.49 159.415 ;
		RECT	2.11 159.285 2.16 159.415 ;
		RECT	3.09 159.285 3.14 159.415 ;
		RECT	4.38 159.285 4.43 159.415 ;
		RECT	6.215 159.285 6.265 159.415 ;
		RECT	3.6 159.055 3.65 159.185 ;
		RECT	1.625 158.595 1.675 158.725 ;
		RECT	1.88 158.635 2.01 158.685 ;
		RECT	5.01 158.635 5.14 158.685 ;
		RECT	3.6 156.635 3.65 156.765 ;
		RECT	1.44 156.405 1.49 156.535 ;
		RECT	2.11 156.405 2.16 156.535 ;
		RECT	3.09 156.405 3.14 156.535 ;
		RECT	4.38 156.405 4.43 156.535 ;
		RECT	6.215 156.405 6.265 156.535 ;
		RECT	3.6 3.535 3.65 3.665 ;
		RECT	1.625 3.075 1.675 3.205 ;
		RECT	1.88 3.115 2.01 3.165 ;
		RECT	5.01 3.115 5.14 3.165 ;
		RECT	3.6 1.115 3.65 1.245 ;
		RECT	1.44 0.885 1.49 1.015 ;
		RECT	2.11 0.885 2.16 1.015 ;
		RECT	3.09 0.885 3.14 1.015 ;
		RECT	4.38 0.885 4.43 1.015 ;
		RECT	6.215 0.885 6.265 1.015 ;
		RECT	3.6 184.975 3.65 185.105 ;
		RECT	1.625 184.515 1.675 184.645 ;
		RECT	1.88 184.555 2.01 184.605 ;
		RECT	5.01 184.555 5.14 184.605 ;
		RECT	3.6 182.555 3.65 182.685 ;
		RECT	1.44 182.325 1.49 182.455 ;
		RECT	2.11 182.325 2.16 182.455 ;
		RECT	3.09 182.325 3.14 182.455 ;
		RECT	4.38 182.325 4.43 182.455 ;
		RECT	6.215 182.325 6.265 182.455 ;
		RECT	0.435 184.515 0.485 184.645 ;
		RECT	0.435 184.975 0.485 185.105 ;
		RECT	0.435 182.555 0.485 182.685 ;
		RECT	0.435 181.635 0.485 181.765 ;
		RECT	0.435 182.095 0.485 182.225 ;
		RECT	0.435 179.675 0.485 179.805 ;
		RECT	0.435 155.715 0.485 155.845 ;
		RECT	0.435 156.175 0.485 156.305 ;
		RECT	0.435 153.755 0.485 153.885 ;
		RECT	0.435 152.835 0.485 152.965 ;
		RECT	0.435 153.295 0.485 153.425 ;
		RECT	0.435 150.875 0.485 151.005 ;
		RECT	0.435 149.955 0.485 150.085 ;
		RECT	0.435 150.415 0.485 150.545 ;
		RECT	0.435 147.995 0.485 148.125 ;
		RECT	0.435 147.075 0.485 147.205 ;
		RECT	0.435 147.535 0.485 147.665 ;
		RECT	0.435 145.115 0.485 145.245 ;
		RECT	0.435 144.195 0.485 144.325 ;
		RECT	0.435 144.655 0.485 144.785 ;
		RECT	0.435 142.235 0.485 142.365 ;
		RECT	0.435 141.315 0.485 141.445 ;
		RECT	0.435 141.775 0.485 141.905 ;
		RECT	0.435 139.355 0.485 139.485 ;
		RECT	0.435 138.435 0.485 138.565 ;
		RECT	0.435 138.895 0.485 139.025 ;
		RECT	0.435 136.475 0.485 136.605 ;
		RECT	0.435 135.555 0.485 135.685 ;
		RECT	0.435 136.015 0.485 136.145 ;
		RECT	0.435 133.595 0.485 133.725 ;
		RECT	0.435 132.675 0.485 132.805 ;
		RECT	0.435 133.135 0.485 133.265 ;
		RECT	0.435 130.715 0.485 130.845 ;
		RECT	0.435 129.795 0.485 129.925 ;
		RECT	0.435 130.255 0.485 130.385 ;
		RECT	0.435 127.835 0.485 127.965 ;
		RECT	0.435 178.755 0.485 178.885 ;
		RECT	0.435 179.215 0.485 179.345 ;
		RECT	0.435 176.795 0.485 176.925 ;
		RECT	0.435 126.915 0.485 127.045 ;
		RECT	0.435 127.375 0.485 127.505 ;
		RECT	0.435 124.955 0.485 125.085 ;
		RECT	0.435 124.035 0.485 124.165 ;
		RECT	0.435 124.495 0.485 124.625 ;
		RECT	0.435 122.075 0.485 122.205 ;
		RECT	0.435 121.155 0.485 121.285 ;
		RECT	0.435 121.615 0.485 121.745 ;
		RECT	0.435 119.195 0.485 119.325 ;
		RECT	0.435 118.275 0.485 118.405 ;
		RECT	0.435 118.735 0.485 118.865 ;
		RECT	0.435 116.315 0.485 116.445 ;
		RECT	0.435 115.395 0.485 115.525 ;
		RECT	0.435 115.855 0.485 115.985 ;
		RECT	0.435 113.435 0.485 113.565 ;
		RECT	0.435 112.515 0.485 112.645 ;
		RECT	0.435 112.975 0.485 113.105 ;
		RECT	0.435 110.555 0.485 110.685 ;
		RECT	0.435 109.635 0.485 109.765 ;
		RECT	0.435 110.095 0.485 110.225 ;
		RECT	0.435 107.675 0.485 107.805 ;
		RECT	0.435 106.755 0.485 106.885 ;
		RECT	0.435 107.215 0.485 107.345 ;
		RECT	0.435 104.795 0.485 104.925 ;
		RECT	0.435 103.875 0.485 104.005 ;
		RECT	0.435 104.335 0.485 104.465 ;
		RECT	0.435 101.915 0.485 102.045 ;
		RECT	0.435 100.995 0.485 101.125 ;
		RECT	0.435 101.455 0.485 101.585 ;
		RECT	0.435 99.035 0.485 99.165 ;
		RECT	0.435 175.875 0.485 176.005 ;
		RECT	0.435 176.335 0.485 176.465 ;
		RECT	0.435 173.915 0.485 174.045 ;
		RECT	0.435 98.115 0.485 98.245 ;
		RECT	0.435 98.575 0.485 98.705 ;
		RECT	0.435 96.155 0.485 96.285 ;
		RECT	0.435 95.235 0.485 95.365 ;
		RECT	0.435 95.695 0.485 95.825 ;
		RECT	0.435 93.275 0.485 93.405 ;
		RECT	0.435 92.355 0.485 92.485 ;
		RECT	0.435 92.815 0.485 92.945 ;
		RECT	0.435 90.395 0.485 90.525 ;
		RECT	0.435 89.475 0.485 89.605 ;
		RECT	0.435 89.935 0.485 90.065 ;
		RECT	0.435 87.515 0.485 87.645 ;
		RECT	0.435 86.595 0.485 86.725 ;
		RECT	0.435 87.055 0.485 87.185 ;
		RECT	0.435 84.635 0.485 84.765 ;
		RECT	0.435 83.715 0.485 83.845 ;
		RECT	0.435 84.175 0.485 84.305 ;
		RECT	0.435 81.755 0.485 81.885 ;
		RECT	0.435 80.835 0.485 80.965 ;
		RECT	0.435 81.295 0.485 81.425 ;
		RECT	0.435 78.875 0.485 79.005 ;
		RECT	0.435 77.955 0.485 78.085 ;
		RECT	0.435 78.415 0.485 78.545 ;
		RECT	0.435 75.995 0.485 76.125 ;
		RECT	0.435 75.075 0.485 75.205 ;
		RECT	0.435 75.535 0.485 75.665 ;
		RECT	0.435 73.115 0.485 73.245 ;
		RECT	0.435 72.195 0.485 72.325 ;
		RECT	0.435 72.655 0.485 72.785 ;
		RECT	0.435 70.235 0.485 70.365 ;
		RECT	0.435 172.995 0.485 173.125 ;
		RECT	0.435 173.455 0.485 173.585 ;
		RECT	0.435 171.035 0.485 171.165 ;
		RECT	0.435 69.315 0.485 69.445 ;
		RECT	0.435 69.775 0.485 69.905 ;
		RECT	0.435 67.355 0.485 67.485 ;
		RECT	0.435 66.435 0.485 66.565 ;
		RECT	0.435 66.895 0.485 67.025 ;
		RECT	0.435 64.475 0.485 64.605 ;
		RECT	0.435 63.555 0.485 63.685 ;
		RECT	0.435 64.015 0.485 64.145 ;
		RECT	0.435 61.595 0.485 61.725 ;
		RECT	0.435 60.675 0.485 60.805 ;
		RECT	0.435 61.135 0.485 61.265 ;
		RECT	0.435 58.715 0.485 58.845 ;
		RECT	0.435 57.795 0.485 57.925 ;
		RECT	0.435 58.255 0.485 58.385 ;
		RECT	0.435 55.835 0.485 55.965 ;
		RECT	0.435 54.915 0.485 55.045 ;
		RECT	0.435 55.375 0.485 55.505 ;
		RECT	0.435 52.955 0.485 53.085 ;
		RECT	0.435 52.035 0.485 52.165 ;
		RECT	0.435 52.495 0.485 52.625 ;
		RECT	0.435 50.075 0.485 50.205 ;
		RECT	0.435 49.155 0.485 49.285 ;
		RECT	0.435 49.615 0.485 49.745 ;
		RECT	0.435 47.195 0.485 47.325 ;
		RECT	0.435 46.275 0.485 46.405 ;
		RECT	0.435 46.735 0.485 46.865 ;
		RECT	0.435 44.315 0.485 44.445 ;
		RECT	0.435 43.395 0.485 43.525 ;
		RECT	0.435 43.855 0.485 43.985 ;
		RECT	0.435 41.435 0.485 41.565 ;
		RECT	0.435 170.115 0.485 170.245 ;
		RECT	0.435 170.575 0.485 170.705 ;
		RECT	0.435 168.155 0.485 168.285 ;
		RECT	0.435 40.515 0.485 40.645 ;
		RECT	0.435 40.975 0.485 41.105 ;
		RECT	0.435 38.555 0.485 38.685 ;
		RECT	0.435 37.635 0.485 37.765 ;
		RECT	0.435 38.095 0.485 38.225 ;
		RECT	0.435 35.675 0.485 35.805 ;
		RECT	0.435 34.755 0.485 34.885 ;
		RECT	0.435 35.215 0.485 35.345 ;
		RECT	0.435 32.795 0.485 32.925 ;
		RECT	0.435 31.875 0.485 32.005 ;
		RECT	0.435 32.335 0.485 32.465 ;
		RECT	0.435 29.915 0.485 30.045 ;
		RECT	0.435 28.995 0.485 29.125 ;
		RECT	0.435 29.455 0.485 29.585 ;
		RECT	0.435 27.035 0.485 27.165 ;
		RECT	0.435 26.115 0.485 26.245 ;
		RECT	0.435 26.575 0.485 26.705 ;
		RECT	0.435 24.155 0.485 24.285 ;
		RECT	0.435 23.235 0.485 23.365 ;
		RECT	0.435 23.695 0.485 23.825 ;
		RECT	0.435 21.275 0.485 21.405 ;
		RECT	0.435 20.355 0.485 20.485 ;
		RECT	0.435 20.815 0.485 20.945 ;
		RECT	0.435 18.395 0.485 18.525 ;
		RECT	0.435 17.475 0.485 17.605 ;
		RECT	0.435 17.935 0.485 18.065 ;
		RECT	0.435 15.515 0.485 15.645 ;
		RECT	0.435 14.595 0.485 14.725 ;
		RECT	0.435 15.055 0.485 15.185 ;
		RECT	0.435 12.635 0.485 12.765 ;
		RECT	0.435 167.235 0.485 167.365 ;
		RECT	0.435 167.695 0.485 167.825 ;
		RECT	0.435 165.275 0.485 165.405 ;
		RECT	0.435 11.715 0.485 11.845 ;
		RECT	0.435 12.175 0.485 12.305 ;
		RECT	0.435 9.755 0.485 9.885 ;
		RECT	0.435 8.835 0.485 8.965 ;
		RECT	0.435 9.295 0.485 9.425 ;
		RECT	0.435 6.875 0.485 7.005 ;
		RECT	0.435 5.955 0.485 6.085 ;
		RECT	0.435 6.415 0.485 6.545 ;
		RECT	0.435 3.995 0.485 4.125 ;
		RECT	0.435 3.075 0.485 3.205 ;
		RECT	0.435 3.535 0.485 3.665 ;
		RECT	0.435 1.115 0.485 1.245 ;
		RECT	0.435 164.355 0.485 164.485 ;
		RECT	0.435 164.815 0.485 164.945 ;
		RECT	0.435 162.395 0.485 162.525 ;
		RECT	0.435 161.475 0.485 161.605 ;
		RECT	0.435 161.935 0.485 162.065 ;
		RECT	0.435 159.515 0.485 159.645 ;
		RECT	0.435 158.595 0.485 158.725 ;
		RECT	0.435 159.055 0.485 159.185 ;
		RECT	0.435 156.635 0.485 156.765 ;
		RECT	6.76 229.755 6.81 229.885 ;
		RECT	8.04 229.755 8.09 229.885 ;
		RECT	9.58 229.755 9.63 229.885 ;
		RECT	9.855 229.755 9.905 229.885 ;
		RECT	10.26 229.755 10.31 229.885 ;
		RECT	11.565 229.755 11.615 229.885 ;
		RECT	13.33 229.755 13.38 229.885 ;
		RECT	6.765 232.175 6.815 232.305 ;
		RECT	8.04 232.175 8.09 232.305 ;
		RECT	9.58 232.175 9.63 232.305 ;
		RECT	9.855 232.175 9.905 232.305 ;
		RECT	11.565 232.175 11.615 232.305 ;
		RECT	13.33 232.175 13.38 232.305 ;
		RECT	7.72 232.405 7.77 232.535 ;
		RECT	14.68 232.405 14.73 232.535 ;
		RECT	9.1 229.755 9.15 229.885 ;
		RECT	10.81 229.755 10.86 229.885 ;
		RECT	9.1 232.175 9.15 232.305 ;
		RECT	10.81 232.175 10.86 232.305 ;
		RECT	6.76 232.635 6.81 232.765 ;
		RECT	8.04 232.635 8.09 232.765 ;
		RECT	9.58 232.635 9.63 232.765 ;
		RECT	9.855 232.635 9.905 232.765 ;
		RECT	10.26 232.635 10.31 232.765 ;
		RECT	11.565 232.635 11.615 232.765 ;
		RECT	13.33 232.635 13.38 232.765 ;
		RECT	6.765 235.055 6.815 235.185 ;
		RECT	8.04 235.055 8.09 235.185 ;
		RECT	9.58 235.055 9.63 235.185 ;
		RECT	9.855 235.055 9.905 235.185 ;
		RECT	11.565 235.055 11.615 235.185 ;
		RECT	13.33 235.055 13.38 235.185 ;
		RECT	7.72 235.285 7.77 235.415 ;
		RECT	14.68 235.285 14.73 235.415 ;
		RECT	9.1 232.635 9.15 232.765 ;
		RECT	10.81 232.635 10.86 232.765 ;
		RECT	9.1 235.055 9.15 235.185 ;
		RECT	10.81 235.055 10.86 235.185 ;
		RECT	6.76 235.515 6.81 235.645 ;
		RECT	8.04 235.515 8.09 235.645 ;
		RECT	9.58 235.515 9.63 235.645 ;
		RECT	9.855 235.515 9.905 235.645 ;
		RECT	10.26 235.515 10.31 235.645 ;
		RECT	11.565 235.515 11.615 235.645 ;
		RECT	13.33 235.515 13.38 235.645 ;
		RECT	6.765 237.935 6.815 238.065 ;
		RECT	8.04 237.935 8.09 238.065 ;
		RECT	9.58 237.935 9.63 238.065 ;
		RECT	9.855 237.935 9.905 238.065 ;
		RECT	11.565 237.935 11.615 238.065 ;
		RECT	13.33 237.935 13.38 238.065 ;
		RECT	7.72 238.165 7.77 238.295 ;
		RECT	14.68 238.165 14.73 238.295 ;
		RECT	9.1 235.515 9.15 235.645 ;
		RECT	10.81 235.515 10.86 235.645 ;
		RECT	9.1 237.935 9.15 238.065 ;
		RECT	10.81 237.935 10.86 238.065 ;
		RECT	6.76 238.395 6.81 238.525 ;
		RECT	8.04 238.395 8.09 238.525 ;
		RECT	9.58 238.395 9.63 238.525 ;
		RECT	9.855 238.395 9.905 238.525 ;
		RECT	10.26 238.395 10.31 238.525 ;
		RECT	11.565 238.395 11.615 238.525 ;
		RECT	13.33 238.395 13.38 238.525 ;
		RECT	6.765 240.815 6.815 240.945 ;
		RECT	8.04 240.815 8.09 240.945 ;
		RECT	9.58 240.815 9.63 240.945 ;
		RECT	9.855 240.815 9.905 240.945 ;
		RECT	11.565 240.815 11.615 240.945 ;
		RECT	13.33 240.815 13.38 240.945 ;
		RECT	7.72 241.045 7.77 241.175 ;
		RECT	14.68 241.045 14.73 241.175 ;
		RECT	9.1 238.395 9.15 238.525 ;
		RECT	10.81 238.395 10.86 238.525 ;
		RECT	9.1 240.815 9.15 240.945 ;
		RECT	10.81 240.815 10.86 240.945 ;
		RECT	6.76 241.275 6.81 241.405 ;
		RECT	8.04 241.275 8.09 241.405 ;
		RECT	9.58 241.275 9.63 241.405 ;
		RECT	9.855 241.275 9.905 241.405 ;
		RECT	10.26 241.275 10.31 241.405 ;
		RECT	11.565 241.275 11.615 241.405 ;
		RECT	13.33 241.275 13.38 241.405 ;
		RECT	6.765 243.695 6.815 243.825 ;
		RECT	8.04 243.695 8.09 243.825 ;
		RECT	9.58 243.695 9.63 243.825 ;
		RECT	9.855 243.695 9.905 243.825 ;
		RECT	11.565 243.695 11.615 243.825 ;
		RECT	13.33 243.695 13.38 243.825 ;
		RECT	7.72 243.925 7.77 244.055 ;
		RECT	14.68 243.925 14.73 244.055 ;
		RECT	9.1 241.275 9.15 241.405 ;
		RECT	10.81 241.275 10.86 241.405 ;
		RECT	9.1 243.695 9.15 243.825 ;
		RECT	10.81 243.695 10.86 243.825 ;
		RECT	6.76 244.155 6.81 244.285 ;
		RECT	8.04 244.155 8.09 244.285 ;
		RECT	9.58 244.155 9.63 244.285 ;
		RECT	9.855 244.155 9.905 244.285 ;
		RECT	10.26 244.155 10.31 244.285 ;
		RECT	11.565 244.155 11.615 244.285 ;
		RECT	13.33 244.155 13.38 244.285 ;
		RECT	6.765 246.575 6.815 246.705 ;
		RECT	8.04 246.575 8.09 246.705 ;
		RECT	9.58 246.575 9.63 246.705 ;
		RECT	9.855 246.575 9.905 246.705 ;
		RECT	11.565 246.575 11.615 246.705 ;
		RECT	13.33 246.575 13.38 246.705 ;
		RECT	7.72 246.805 7.77 246.935 ;
		RECT	14.68 246.805 14.73 246.935 ;
		RECT	9.1 244.155 9.15 244.285 ;
		RECT	10.81 244.155 10.86 244.285 ;
		RECT	9.1 246.575 9.15 246.705 ;
		RECT	10.81 246.575 10.86 246.705 ;
		RECT	6.76 247.035 6.81 247.165 ;
		RECT	8.04 247.035 8.09 247.165 ;
		RECT	9.58 247.035 9.63 247.165 ;
		RECT	9.855 247.035 9.905 247.165 ;
		RECT	10.26 247.035 10.31 247.165 ;
		RECT	11.565 247.035 11.615 247.165 ;
		RECT	13.33 247.035 13.38 247.165 ;
		RECT	6.765 249.455 6.815 249.585 ;
		RECT	8.04 249.455 8.09 249.585 ;
		RECT	9.58 249.455 9.63 249.585 ;
		RECT	9.855 249.455 9.905 249.585 ;
		RECT	11.565 249.455 11.615 249.585 ;
		RECT	13.33 249.455 13.38 249.585 ;
		RECT	7.72 249.685 7.77 249.815 ;
		RECT	14.68 249.685 14.73 249.815 ;
		RECT	9.1 247.035 9.15 247.165 ;
		RECT	10.81 247.035 10.86 247.165 ;
		RECT	9.1 249.455 9.15 249.585 ;
		RECT	10.81 249.455 10.86 249.585 ;
		RECT	6.76 249.915 6.81 250.045 ;
		RECT	8.04 249.915 8.09 250.045 ;
		RECT	9.58 249.915 9.63 250.045 ;
		RECT	9.855 249.915 9.905 250.045 ;
		RECT	10.26 249.915 10.31 250.045 ;
		RECT	11.565 249.915 11.615 250.045 ;
		RECT	13.33 249.915 13.38 250.045 ;
		RECT	6.765 252.335 6.815 252.465 ;
		RECT	8.04 252.335 8.09 252.465 ;
		RECT	9.58 252.335 9.63 252.465 ;
		RECT	9.855 252.335 9.905 252.465 ;
		RECT	11.565 252.335 11.615 252.465 ;
		RECT	13.33 252.335 13.38 252.465 ;
		RECT	7.72 252.565 7.77 252.695 ;
		RECT	14.68 252.565 14.73 252.695 ;
		RECT	9.1 249.915 9.15 250.045 ;
		RECT	10.81 249.915 10.86 250.045 ;
		RECT	9.1 252.335 9.15 252.465 ;
		RECT	10.81 252.335 10.86 252.465 ;
		RECT	6.76 252.795 6.81 252.925 ;
		RECT	8.04 252.795 8.09 252.925 ;
		RECT	9.58 252.795 9.63 252.925 ;
		RECT	9.855 252.795 9.905 252.925 ;
		RECT	10.26 252.795 10.31 252.925 ;
		RECT	11.565 252.795 11.615 252.925 ;
		RECT	13.33 252.795 13.38 252.925 ;
		RECT	6.765 255.215 6.815 255.345 ;
		RECT	8.04 255.215 8.09 255.345 ;
		RECT	9.58 255.215 9.63 255.345 ;
		RECT	9.855 255.215 9.905 255.345 ;
		RECT	11.565 255.215 11.615 255.345 ;
		RECT	13.33 255.215 13.38 255.345 ;
		RECT	7.72 255.445 7.77 255.575 ;
		RECT	14.68 255.445 14.73 255.575 ;
		RECT	9.1 252.795 9.15 252.925 ;
		RECT	10.81 252.795 10.86 252.925 ;
		RECT	9.1 255.215 9.15 255.345 ;
		RECT	10.81 255.215 10.86 255.345 ;
		RECT	6.76 255.675 6.81 255.805 ;
		RECT	8.04 255.675 8.09 255.805 ;
		RECT	9.58 255.675 9.63 255.805 ;
		RECT	9.855 255.675 9.905 255.805 ;
		RECT	10.26 255.675 10.31 255.805 ;
		RECT	11.565 255.675 11.615 255.805 ;
		RECT	13.33 255.675 13.38 255.805 ;
		RECT	6.765 258.095 6.815 258.225 ;
		RECT	8.04 258.095 8.09 258.225 ;
		RECT	9.58 258.095 9.63 258.225 ;
		RECT	9.855 258.095 9.905 258.225 ;
		RECT	11.565 258.095 11.615 258.225 ;
		RECT	13.33 258.095 13.38 258.225 ;
		RECT	7.72 258.325 7.77 258.455 ;
		RECT	14.68 258.325 14.73 258.455 ;
		RECT	9.1 255.675 9.15 255.805 ;
		RECT	10.81 255.675 10.86 255.805 ;
		RECT	9.1 258.095 9.15 258.225 ;
		RECT	10.81 258.095 10.86 258.225 ;
		RECT	6.76 258.555 6.81 258.685 ;
		RECT	8.04 258.555 8.09 258.685 ;
		RECT	9.58 258.555 9.63 258.685 ;
		RECT	9.855 258.555 9.905 258.685 ;
		RECT	10.26 258.555 10.31 258.685 ;
		RECT	11.565 258.555 11.615 258.685 ;
		RECT	13.33 258.555 13.38 258.685 ;
		RECT	6.765 260.975 6.815 261.105 ;
		RECT	8.04 260.975 8.09 261.105 ;
		RECT	9.58 260.975 9.63 261.105 ;
		RECT	9.855 260.975 9.905 261.105 ;
		RECT	11.565 260.975 11.615 261.105 ;
		RECT	13.33 260.975 13.38 261.105 ;
		RECT	7.72 261.205 7.77 261.335 ;
		RECT	14.68 261.205 14.73 261.335 ;
		RECT	9.1 258.555 9.15 258.685 ;
		RECT	10.81 258.555 10.86 258.685 ;
		RECT	9.1 260.975 9.15 261.105 ;
		RECT	10.81 260.975 10.86 261.105 ;
		RECT	6.76 261.435 6.81 261.565 ;
		RECT	8.04 261.435 8.09 261.565 ;
		RECT	9.58 261.435 9.63 261.565 ;
		RECT	9.855 261.435 9.905 261.565 ;
		RECT	10.26 261.435 10.31 261.565 ;
		RECT	11.565 261.435 11.615 261.565 ;
		RECT	13.33 261.435 13.38 261.565 ;
		RECT	6.765 263.855 6.815 263.985 ;
		RECT	8.04 263.855 8.09 263.985 ;
		RECT	9.58 263.855 9.63 263.985 ;
		RECT	9.855 263.855 9.905 263.985 ;
		RECT	11.565 263.855 11.615 263.985 ;
		RECT	13.33 263.855 13.38 263.985 ;
		RECT	7.72 264.085 7.77 264.215 ;
		RECT	14.68 264.085 14.73 264.215 ;
		RECT	9.1 261.435 9.15 261.565 ;
		RECT	10.81 261.435 10.86 261.565 ;
		RECT	9.1 263.855 9.15 263.985 ;
		RECT	10.81 263.855 10.86 263.985 ;
		RECT	6.76 264.315 6.81 264.445 ;
		RECT	8.04 264.315 8.09 264.445 ;
		RECT	9.58 264.315 9.63 264.445 ;
		RECT	9.855 264.315 9.905 264.445 ;
		RECT	10.26 264.315 10.31 264.445 ;
		RECT	11.565 264.315 11.615 264.445 ;
		RECT	13.33 264.315 13.38 264.445 ;
		RECT	6.765 266.735 6.815 266.865 ;
		RECT	8.04 266.735 8.09 266.865 ;
		RECT	9.58 266.735 9.63 266.865 ;
		RECT	9.855 266.735 9.905 266.865 ;
		RECT	11.565 266.735 11.615 266.865 ;
		RECT	13.33 266.735 13.38 266.865 ;
		RECT	7.72 266.965 7.77 267.095 ;
		RECT	14.68 266.965 14.73 267.095 ;
		RECT	9.1 264.315 9.15 264.445 ;
		RECT	10.81 264.315 10.86 264.445 ;
		RECT	9.1 266.735 9.15 266.865 ;
		RECT	10.81 266.735 10.86 266.865 ;
		RECT	6.76 267.195 6.81 267.325 ;
		RECT	8.04 267.195 8.09 267.325 ;
		RECT	9.58 267.195 9.63 267.325 ;
		RECT	9.855 267.195 9.905 267.325 ;
		RECT	10.26 267.195 10.31 267.325 ;
		RECT	11.565 267.195 11.615 267.325 ;
		RECT	13.33 267.195 13.38 267.325 ;
		RECT	6.765 269.615 6.815 269.745 ;
		RECT	8.04 269.615 8.09 269.745 ;
		RECT	9.58 269.615 9.63 269.745 ;
		RECT	9.855 269.615 9.905 269.745 ;
		RECT	11.565 269.615 11.615 269.745 ;
		RECT	13.33 269.615 13.38 269.745 ;
		RECT	7.72 269.845 7.77 269.975 ;
		RECT	14.68 269.845 14.73 269.975 ;
		RECT	9.1 267.195 9.15 267.325 ;
		RECT	10.81 267.195 10.86 267.325 ;
		RECT	9.1 269.615 9.15 269.745 ;
		RECT	10.81 269.615 10.86 269.745 ;
		RECT	6.76 270.075 6.81 270.205 ;
		RECT	8.04 270.075 8.09 270.205 ;
		RECT	9.58 270.075 9.63 270.205 ;
		RECT	9.855 270.075 9.905 270.205 ;
		RECT	10.26 270.075 10.31 270.205 ;
		RECT	11.565 270.075 11.615 270.205 ;
		RECT	13.33 270.075 13.38 270.205 ;
		RECT	6.765 272.495 6.815 272.625 ;
		RECT	8.04 272.495 8.09 272.625 ;
		RECT	9.58 272.495 9.63 272.625 ;
		RECT	9.855 272.495 9.905 272.625 ;
		RECT	11.565 272.495 11.615 272.625 ;
		RECT	13.33 272.495 13.38 272.625 ;
		RECT	7.72 272.725 7.77 272.855 ;
		RECT	14.68 272.725 14.73 272.855 ;
		RECT	9.1 270.075 9.15 270.205 ;
		RECT	10.81 270.075 10.86 270.205 ;
		RECT	9.1 272.495 9.15 272.625 ;
		RECT	10.81 272.495 10.86 272.625 ;
		RECT	6.76 272.955 6.81 273.085 ;
		RECT	8.04 272.955 8.09 273.085 ;
		RECT	9.58 272.955 9.63 273.085 ;
		RECT	9.855 272.955 9.905 273.085 ;
		RECT	10.26 272.955 10.31 273.085 ;
		RECT	11.565 272.955 11.615 273.085 ;
		RECT	13.33 272.955 13.38 273.085 ;
		RECT	6.765 275.375 6.815 275.505 ;
		RECT	8.04 275.375 8.09 275.505 ;
		RECT	9.58 275.375 9.63 275.505 ;
		RECT	9.855 275.375 9.905 275.505 ;
		RECT	11.565 275.375 11.615 275.505 ;
		RECT	13.33 275.375 13.38 275.505 ;
		RECT	7.72 275.605 7.77 275.735 ;
		RECT	14.68 275.605 14.73 275.735 ;
		RECT	9.1 272.955 9.15 273.085 ;
		RECT	10.81 272.955 10.86 273.085 ;
		RECT	9.1 275.375 9.15 275.505 ;
		RECT	10.81 275.375 10.86 275.505 ;
		RECT	6.76 275.835 6.81 275.965 ;
		RECT	8.04 275.835 8.09 275.965 ;
		RECT	9.58 275.835 9.63 275.965 ;
		RECT	9.855 275.835 9.905 275.965 ;
		RECT	10.26 275.835 10.31 275.965 ;
		RECT	11.565 275.835 11.615 275.965 ;
		RECT	13.33 275.835 13.38 275.965 ;
		RECT	6.765 278.255 6.815 278.385 ;
		RECT	8.04 278.255 8.09 278.385 ;
		RECT	9.58 278.255 9.63 278.385 ;
		RECT	9.855 278.255 9.905 278.385 ;
		RECT	11.565 278.255 11.615 278.385 ;
		RECT	13.33 278.255 13.38 278.385 ;
		RECT	7.72 278.485 7.77 278.615 ;
		RECT	14.68 278.485 14.73 278.615 ;
		RECT	9.1 275.835 9.15 275.965 ;
		RECT	10.81 275.835 10.86 275.965 ;
		RECT	9.1 278.255 9.15 278.385 ;
		RECT	10.81 278.255 10.86 278.385 ;
		RECT	6.76 278.715 6.81 278.845 ;
		RECT	8.04 278.715 8.09 278.845 ;
		RECT	9.58 278.715 9.63 278.845 ;
		RECT	9.855 278.715 9.905 278.845 ;
		RECT	10.26 278.715 10.31 278.845 ;
		RECT	11.565 278.715 11.615 278.845 ;
		RECT	13.33 278.715 13.38 278.845 ;
		RECT	6.765 281.135 6.815 281.265 ;
		RECT	8.04 281.135 8.09 281.265 ;
		RECT	9.58 281.135 9.63 281.265 ;
		RECT	9.855 281.135 9.905 281.265 ;
		RECT	11.565 281.135 11.615 281.265 ;
		RECT	13.33 281.135 13.38 281.265 ;
		RECT	7.72 281.365 7.77 281.495 ;
		RECT	14.68 281.365 14.73 281.495 ;
		RECT	9.1 278.715 9.15 278.845 ;
		RECT	10.81 278.715 10.86 278.845 ;
		RECT	9.1 281.135 9.15 281.265 ;
		RECT	10.81 281.135 10.86 281.265 ;
		RECT	6.76 281.595 6.81 281.725 ;
		RECT	8.04 281.595 8.09 281.725 ;
		RECT	9.58 281.595 9.63 281.725 ;
		RECT	9.855 281.595 9.905 281.725 ;
		RECT	10.26 281.595 10.31 281.725 ;
		RECT	11.565 281.595 11.615 281.725 ;
		RECT	13.33 281.595 13.38 281.725 ;
		RECT	6.765 284.015 6.815 284.145 ;
		RECT	8.04 284.015 8.09 284.145 ;
		RECT	9.58 284.015 9.63 284.145 ;
		RECT	9.855 284.015 9.905 284.145 ;
		RECT	11.565 284.015 11.615 284.145 ;
		RECT	13.33 284.015 13.38 284.145 ;
		RECT	7.72 284.245 7.77 284.375 ;
		RECT	14.68 284.245 14.73 284.375 ;
		RECT	9.1 281.595 9.15 281.725 ;
		RECT	10.81 281.595 10.86 281.725 ;
		RECT	9.1 284.015 9.15 284.145 ;
		RECT	10.81 284.015 10.86 284.145 ;
		RECT	6.76 284.475 6.81 284.605 ;
		RECT	8.04 284.475 8.09 284.605 ;
		RECT	9.58 284.475 9.63 284.605 ;
		RECT	9.855 284.475 9.905 284.605 ;
		RECT	10.26 284.475 10.31 284.605 ;
		RECT	11.565 284.475 11.615 284.605 ;
		RECT	13.33 284.475 13.38 284.605 ;
		RECT	6.765 286.895 6.815 287.025 ;
		RECT	8.04 286.895 8.09 287.025 ;
		RECT	9.58 286.895 9.63 287.025 ;
		RECT	9.855 286.895 9.905 287.025 ;
		RECT	11.565 286.895 11.615 287.025 ;
		RECT	13.33 286.895 13.38 287.025 ;
		RECT	7.72 287.125 7.77 287.255 ;
		RECT	14.68 287.125 14.73 287.255 ;
		RECT	9.1 284.475 9.15 284.605 ;
		RECT	10.81 284.475 10.86 284.605 ;
		RECT	9.1 286.895 9.15 287.025 ;
		RECT	10.81 286.895 10.86 287.025 ;
		RECT	6.76 287.355 6.81 287.485 ;
		RECT	8.04 287.355 8.09 287.485 ;
		RECT	9.58 287.355 9.63 287.485 ;
		RECT	9.855 287.355 9.905 287.485 ;
		RECT	10.26 287.355 10.31 287.485 ;
		RECT	11.565 287.355 11.615 287.485 ;
		RECT	13.33 287.355 13.38 287.485 ;
		RECT	6.765 289.775 6.815 289.905 ;
		RECT	8.04 289.775 8.09 289.905 ;
		RECT	9.58 289.775 9.63 289.905 ;
		RECT	9.855 289.775 9.905 289.905 ;
		RECT	11.565 289.775 11.615 289.905 ;
		RECT	13.33 289.775 13.38 289.905 ;
		RECT	7.72 290.005 7.77 290.135 ;
		RECT	14.68 290.005 14.73 290.135 ;
		RECT	9.1 287.355 9.15 287.485 ;
		RECT	10.81 287.355 10.86 287.485 ;
		RECT	9.1 289.775 9.15 289.905 ;
		RECT	10.81 289.775 10.86 289.905 ;
		RECT	6.76 290.235 6.81 290.365 ;
		RECT	8.04 290.235 8.09 290.365 ;
		RECT	9.58 290.235 9.63 290.365 ;
		RECT	9.855 290.235 9.905 290.365 ;
		RECT	10.26 290.235 10.31 290.365 ;
		RECT	11.565 290.235 11.615 290.365 ;
		RECT	13.33 290.235 13.38 290.365 ;
		RECT	6.765 292.655 6.815 292.785 ;
		RECT	8.04 292.655 8.09 292.785 ;
		RECT	9.58 292.655 9.63 292.785 ;
		RECT	9.855 292.655 9.905 292.785 ;
		RECT	11.565 292.655 11.615 292.785 ;
		RECT	13.33 292.655 13.38 292.785 ;
		RECT	7.72 292.885 7.77 293.015 ;
		RECT	14.68 292.885 14.73 293.015 ;
		RECT	9.1 290.235 9.15 290.365 ;
		RECT	10.81 290.235 10.86 290.365 ;
		RECT	9.1 292.655 9.15 292.785 ;
		RECT	10.81 292.655 10.86 292.785 ;
		RECT	6.76 293.115 6.81 293.245 ;
		RECT	8.04 293.115 8.09 293.245 ;
		RECT	9.58 293.115 9.63 293.245 ;
		RECT	9.855 293.115 9.905 293.245 ;
		RECT	10.26 293.115 10.31 293.245 ;
		RECT	11.565 293.115 11.615 293.245 ;
		RECT	13.33 293.115 13.38 293.245 ;
		RECT	6.765 295.535 6.815 295.665 ;
		RECT	8.04 295.535 8.09 295.665 ;
		RECT	9.58 295.535 9.63 295.665 ;
		RECT	9.855 295.535 9.905 295.665 ;
		RECT	11.565 295.535 11.615 295.665 ;
		RECT	13.33 295.535 13.38 295.665 ;
		RECT	7.72 295.765 7.77 295.895 ;
		RECT	14.68 295.765 14.73 295.895 ;
		RECT	9.1 293.115 9.15 293.245 ;
		RECT	10.81 293.115 10.86 293.245 ;
		RECT	9.1 295.535 9.15 295.665 ;
		RECT	10.81 295.535 10.86 295.665 ;
		RECT	6.76 295.995 6.81 296.125 ;
		RECT	8.04 295.995 8.09 296.125 ;
		RECT	9.58 295.995 9.63 296.125 ;
		RECT	9.855 295.995 9.905 296.125 ;
		RECT	10.26 295.995 10.31 296.125 ;
		RECT	11.565 295.995 11.615 296.125 ;
		RECT	13.33 295.995 13.38 296.125 ;
		RECT	6.765 298.415 6.815 298.545 ;
		RECT	8.04 298.415 8.09 298.545 ;
		RECT	9.58 298.415 9.63 298.545 ;
		RECT	9.855 298.415 9.905 298.545 ;
		RECT	11.565 298.415 11.615 298.545 ;
		RECT	13.33 298.415 13.38 298.545 ;
		RECT	7.72 298.645 7.77 298.775 ;
		RECT	14.68 298.645 14.73 298.775 ;
		RECT	9.1 295.995 9.15 296.125 ;
		RECT	10.81 295.995 10.86 296.125 ;
		RECT	9.1 298.415 9.15 298.545 ;
		RECT	10.81 298.415 10.86 298.545 ;
		RECT	6.76 298.875 6.81 299.005 ;
		RECT	8.04 298.875 8.09 299.005 ;
		RECT	9.58 298.875 9.63 299.005 ;
		RECT	9.855 298.875 9.905 299.005 ;
		RECT	10.26 298.875 10.31 299.005 ;
		RECT	11.565 298.875 11.615 299.005 ;
		RECT	13.33 298.875 13.38 299.005 ;
		RECT	6.765 301.295 6.815 301.425 ;
		RECT	8.04 301.295 8.09 301.425 ;
		RECT	9.58 301.295 9.63 301.425 ;
		RECT	9.855 301.295 9.905 301.425 ;
		RECT	11.565 301.295 11.615 301.425 ;
		RECT	13.33 301.295 13.38 301.425 ;
		RECT	7.72 301.525 7.77 301.655 ;
		RECT	14.68 301.525 14.73 301.655 ;
		RECT	9.1 298.875 9.15 299.005 ;
		RECT	10.81 298.875 10.86 299.005 ;
		RECT	9.1 301.295 9.15 301.425 ;
		RECT	10.81 301.295 10.86 301.425 ;
		RECT	6.76 301.755 6.81 301.885 ;
		RECT	8.04 301.755 8.09 301.885 ;
		RECT	9.58 301.755 9.63 301.885 ;
		RECT	9.855 301.755 9.905 301.885 ;
		RECT	10.26 301.755 10.31 301.885 ;
		RECT	11.565 301.755 11.615 301.885 ;
		RECT	13.33 301.755 13.38 301.885 ;
		RECT	6.765 304.175 6.815 304.305 ;
		RECT	8.04 304.175 8.09 304.305 ;
		RECT	9.58 304.175 9.63 304.305 ;
		RECT	9.855 304.175 9.905 304.305 ;
		RECT	11.565 304.175 11.615 304.305 ;
		RECT	13.33 304.175 13.38 304.305 ;
		RECT	7.72 304.405 7.77 304.535 ;
		RECT	14.68 304.405 14.73 304.535 ;
		RECT	9.1 301.755 9.15 301.885 ;
		RECT	10.81 301.755 10.86 301.885 ;
		RECT	9.1 304.175 9.15 304.305 ;
		RECT	10.81 304.175 10.86 304.305 ;
		RECT	6.76 304.635 6.81 304.765 ;
		RECT	8.04 304.635 8.09 304.765 ;
		RECT	9.58 304.635 9.63 304.765 ;
		RECT	9.855 304.635 9.905 304.765 ;
		RECT	10.26 304.635 10.31 304.765 ;
		RECT	11.565 304.635 11.615 304.765 ;
		RECT	13.33 304.635 13.38 304.765 ;
		RECT	6.765 307.055 6.815 307.185 ;
		RECT	8.04 307.055 8.09 307.185 ;
		RECT	9.58 307.055 9.63 307.185 ;
		RECT	9.855 307.055 9.905 307.185 ;
		RECT	11.565 307.055 11.615 307.185 ;
		RECT	13.33 307.055 13.38 307.185 ;
		RECT	7.72 307.285 7.77 307.415 ;
		RECT	14.68 307.285 14.73 307.415 ;
		RECT	9.1 304.635 9.15 304.765 ;
		RECT	10.81 304.635 10.86 304.765 ;
		RECT	9.1 307.055 9.15 307.185 ;
		RECT	10.81 307.055 10.86 307.185 ;
		RECT	6.76 307.515 6.81 307.645 ;
		RECT	8.04 307.515 8.09 307.645 ;
		RECT	9.58 307.515 9.63 307.645 ;
		RECT	9.855 307.515 9.905 307.645 ;
		RECT	10.26 307.515 10.31 307.645 ;
		RECT	11.565 307.515 11.615 307.645 ;
		RECT	13.33 307.515 13.38 307.645 ;
		RECT	6.765 309.935 6.815 310.065 ;
		RECT	8.04 309.935 8.09 310.065 ;
		RECT	9.58 309.935 9.63 310.065 ;
		RECT	9.855 309.935 9.905 310.065 ;
		RECT	11.565 309.935 11.615 310.065 ;
		RECT	13.33 309.935 13.38 310.065 ;
		RECT	7.72 310.165 7.77 310.295 ;
		RECT	14.68 310.165 14.73 310.295 ;
		RECT	9.1 307.515 9.15 307.645 ;
		RECT	10.81 307.515 10.86 307.645 ;
		RECT	9.1 309.935 9.15 310.065 ;
		RECT	10.81 309.935 10.86 310.065 ;
		RECT	6.76 310.395 6.81 310.525 ;
		RECT	8.04 310.395 8.09 310.525 ;
		RECT	9.58 310.395 9.63 310.525 ;
		RECT	9.855 310.395 9.905 310.525 ;
		RECT	10.26 310.395 10.31 310.525 ;
		RECT	11.565 310.395 11.615 310.525 ;
		RECT	13.33 310.395 13.38 310.525 ;
		RECT	6.765 312.815 6.815 312.945 ;
		RECT	8.04 312.815 8.09 312.945 ;
		RECT	9.58 312.815 9.63 312.945 ;
		RECT	9.855 312.815 9.905 312.945 ;
		RECT	11.565 312.815 11.615 312.945 ;
		RECT	13.33 312.815 13.38 312.945 ;
		RECT	7.72 313.045 7.77 313.175 ;
		RECT	14.68 313.045 14.73 313.175 ;
		RECT	9.1 310.395 9.15 310.525 ;
		RECT	10.81 310.395 10.86 310.525 ;
		RECT	9.1 312.815 9.15 312.945 ;
		RECT	10.81 312.815 10.86 312.945 ;
		RECT	6.76 313.275 6.81 313.405 ;
		RECT	8.04 313.275 8.09 313.405 ;
		RECT	9.58 313.275 9.63 313.405 ;
		RECT	9.855 313.275 9.905 313.405 ;
		RECT	10.26 313.275 10.31 313.405 ;
		RECT	11.565 313.275 11.615 313.405 ;
		RECT	13.33 313.275 13.38 313.405 ;
		RECT	6.765 315.695 6.815 315.825 ;
		RECT	8.04 315.695 8.09 315.825 ;
		RECT	9.58 315.695 9.63 315.825 ;
		RECT	9.855 315.695 9.905 315.825 ;
		RECT	11.565 315.695 11.615 315.825 ;
		RECT	13.33 315.695 13.38 315.825 ;
		RECT	7.72 315.925 7.77 316.055 ;
		RECT	14.68 315.925 14.73 316.055 ;
		RECT	9.1 313.275 9.15 313.405 ;
		RECT	10.81 313.275 10.86 313.405 ;
		RECT	9.1 315.695 9.15 315.825 ;
		RECT	10.81 315.695 10.86 315.825 ;
		RECT	6.76 316.155 6.81 316.285 ;
		RECT	8.04 316.155 8.09 316.285 ;
		RECT	9.58 316.155 9.63 316.285 ;
		RECT	9.855 316.155 9.905 316.285 ;
		RECT	10.26 316.155 10.31 316.285 ;
		RECT	11.565 316.155 11.615 316.285 ;
		RECT	13.33 316.155 13.38 316.285 ;
		RECT	6.765 318.575 6.815 318.705 ;
		RECT	8.04 318.575 8.09 318.705 ;
		RECT	9.58 318.575 9.63 318.705 ;
		RECT	9.855 318.575 9.905 318.705 ;
		RECT	11.565 318.575 11.615 318.705 ;
		RECT	13.33 318.575 13.38 318.705 ;
		RECT	7.72 318.805 7.77 318.935 ;
		RECT	14.68 318.805 14.73 318.935 ;
		RECT	9.1 316.155 9.15 316.285 ;
		RECT	10.81 316.155 10.86 316.285 ;
		RECT	9.1 318.575 9.15 318.705 ;
		RECT	10.81 318.575 10.86 318.705 ;
		RECT	6.76 319.035 6.81 319.165 ;
		RECT	8.04 319.035 8.09 319.165 ;
		RECT	9.58 319.035 9.63 319.165 ;
		RECT	9.855 319.035 9.905 319.165 ;
		RECT	10.26 319.035 10.31 319.165 ;
		RECT	11.565 319.035 11.615 319.165 ;
		RECT	13.33 319.035 13.38 319.165 ;
		RECT	6.765 321.455 6.815 321.585 ;
		RECT	8.04 321.455 8.09 321.585 ;
		RECT	9.58 321.455 9.63 321.585 ;
		RECT	9.855 321.455 9.905 321.585 ;
		RECT	11.565 321.455 11.615 321.585 ;
		RECT	13.33 321.455 13.38 321.585 ;
		RECT	7.72 321.685 7.77 321.815 ;
		RECT	14.68 321.685 14.73 321.815 ;
		RECT	9.1 319.035 9.15 319.165 ;
		RECT	10.81 319.035 10.86 319.165 ;
		RECT	9.1 321.455 9.15 321.585 ;
		RECT	10.81 321.455 10.86 321.585 ;
		RECT	6.76 321.915 6.81 322.045 ;
		RECT	8.04 321.915 8.09 322.045 ;
		RECT	9.58 321.915 9.63 322.045 ;
		RECT	9.855 321.915 9.905 322.045 ;
		RECT	10.26 321.915 10.31 322.045 ;
		RECT	11.565 321.915 11.615 322.045 ;
		RECT	13.33 321.915 13.38 322.045 ;
		RECT	6.765 324.335 6.815 324.465 ;
		RECT	8.04 324.335 8.09 324.465 ;
		RECT	9.58 324.335 9.63 324.465 ;
		RECT	9.855 324.335 9.905 324.465 ;
		RECT	11.565 324.335 11.615 324.465 ;
		RECT	13.33 324.335 13.38 324.465 ;
		RECT	7.72 324.565 7.77 324.695 ;
		RECT	14.68 324.565 14.73 324.695 ;
		RECT	9.1 321.915 9.15 322.045 ;
		RECT	10.81 321.915 10.86 322.045 ;
		RECT	9.1 324.335 9.15 324.465 ;
		RECT	10.81 324.335 10.86 324.465 ;
		RECT	6.76 324.795 6.81 324.925 ;
		RECT	8.04 324.795 8.09 324.925 ;
		RECT	9.58 324.795 9.63 324.925 ;
		RECT	9.855 324.795 9.905 324.925 ;
		RECT	10.26 324.795 10.31 324.925 ;
		RECT	11.565 324.795 11.615 324.925 ;
		RECT	13.33 324.795 13.38 324.925 ;
		RECT	6.765 327.215 6.815 327.345 ;
		RECT	8.04 327.215 8.09 327.345 ;
		RECT	9.58 327.215 9.63 327.345 ;
		RECT	9.855 327.215 9.905 327.345 ;
		RECT	11.565 327.215 11.615 327.345 ;
		RECT	13.33 327.215 13.38 327.345 ;
		RECT	7.72 327.445 7.77 327.575 ;
		RECT	14.68 327.445 14.73 327.575 ;
		RECT	9.1 324.795 9.15 324.925 ;
		RECT	10.81 324.795 10.86 324.925 ;
		RECT	9.1 327.215 9.15 327.345 ;
		RECT	10.81 327.215 10.86 327.345 ;
		RECT	6.76 327.675 6.81 327.805 ;
		RECT	8.04 327.675 8.09 327.805 ;
		RECT	9.58 327.675 9.63 327.805 ;
		RECT	9.855 327.675 9.905 327.805 ;
		RECT	10.26 327.675 10.31 327.805 ;
		RECT	11.565 327.675 11.615 327.805 ;
		RECT	13.33 327.675 13.38 327.805 ;
		RECT	6.765 330.095 6.815 330.225 ;
		RECT	8.04 330.095 8.09 330.225 ;
		RECT	9.58 330.095 9.63 330.225 ;
		RECT	9.855 330.095 9.905 330.225 ;
		RECT	11.565 330.095 11.615 330.225 ;
		RECT	13.33 330.095 13.38 330.225 ;
		RECT	7.72 330.325 7.77 330.455 ;
		RECT	14.68 330.325 14.73 330.455 ;
		RECT	9.1 327.675 9.15 327.805 ;
		RECT	10.81 327.675 10.86 327.805 ;
		RECT	9.1 330.095 9.15 330.225 ;
		RECT	10.81 330.095 10.86 330.225 ;
		RECT	6.76 330.555 6.81 330.685 ;
		RECT	8.04 330.555 8.09 330.685 ;
		RECT	9.58 330.555 9.63 330.685 ;
		RECT	9.855 330.555 9.905 330.685 ;
		RECT	10.26 330.555 10.31 330.685 ;
		RECT	11.565 330.555 11.615 330.685 ;
		RECT	13.33 330.555 13.38 330.685 ;
		RECT	6.765 332.975 6.815 333.105 ;
		RECT	8.04 332.975 8.09 333.105 ;
		RECT	9.58 332.975 9.63 333.105 ;
		RECT	9.855 332.975 9.905 333.105 ;
		RECT	11.565 332.975 11.615 333.105 ;
		RECT	13.33 332.975 13.38 333.105 ;
		RECT	7.72 333.205 7.77 333.335 ;
		RECT	14.68 333.205 14.73 333.335 ;
		RECT	9.1 330.555 9.15 330.685 ;
		RECT	10.81 330.555 10.86 330.685 ;
		RECT	9.1 332.975 9.15 333.105 ;
		RECT	10.81 332.975 10.86 333.105 ;
		RECT	6.76 333.435 6.81 333.565 ;
		RECT	8.04 333.435 8.09 333.565 ;
		RECT	9.58 333.435 9.63 333.565 ;
		RECT	9.855 333.435 9.905 333.565 ;
		RECT	10.26 333.435 10.31 333.565 ;
		RECT	11.565 333.435 11.615 333.565 ;
		RECT	13.33 333.435 13.38 333.565 ;
		RECT	6.765 335.855 6.815 335.985 ;
		RECT	8.04 335.855 8.09 335.985 ;
		RECT	9.58 335.855 9.63 335.985 ;
		RECT	9.855 335.855 9.905 335.985 ;
		RECT	11.565 335.855 11.615 335.985 ;
		RECT	13.33 335.855 13.38 335.985 ;
		RECT	7.72 336.085 7.77 336.215 ;
		RECT	14.68 336.085 14.73 336.215 ;
		RECT	9.1 333.435 9.15 333.565 ;
		RECT	10.81 333.435 10.86 333.565 ;
		RECT	9.1 335.855 9.15 335.985 ;
		RECT	10.81 335.855 10.86 335.985 ;
		RECT	6.76 336.315 6.81 336.445 ;
		RECT	8.04 336.315 8.09 336.445 ;
		RECT	9.58 336.315 9.63 336.445 ;
		RECT	9.855 336.315 9.905 336.445 ;
		RECT	10.26 336.315 10.31 336.445 ;
		RECT	11.565 336.315 11.615 336.445 ;
		RECT	13.33 336.315 13.38 336.445 ;
		RECT	6.765 338.735 6.815 338.865 ;
		RECT	8.04 338.735 8.09 338.865 ;
		RECT	9.58 338.735 9.63 338.865 ;
		RECT	9.855 338.735 9.905 338.865 ;
		RECT	11.565 338.735 11.615 338.865 ;
		RECT	13.33 338.735 13.38 338.865 ;
		RECT	7.72 338.965 7.77 339.095 ;
		RECT	14.68 338.965 14.73 339.095 ;
		RECT	9.1 336.315 9.15 336.445 ;
		RECT	10.81 336.315 10.86 336.445 ;
		RECT	9.1 338.735 9.15 338.865 ;
		RECT	10.81 338.735 10.86 338.865 ;
		RECT	6.76 339.195 6.81 339.325 ;
		RECT	8.04 339.195 8.09 339.325 ;
		RECT	9.58 339.195 9.63 339.325 ;
		RECT	9.855 339.195 9.905 339.325 ;
		RECT	10.26 339.195 10.31 339.325 ;
		RECT	11.565 339.195 11.615 339.325 ;
		RECT	13.33 339.195 13.38 339.325 ;
		RECT	6.765 341.615 6.815 341.745 ;
		RECT	8.04 341.615 8.09 341.745 ;
		RECT	9.58 341.615 9.63 341.745 ;
		RECT	9.855 341.615 9.905 341.745 ;
		RECT	11.565 341.615 11.615 341.745 ;
		RECT	13.33 341.615 13.38 341.745 ;
		RECT	7.72 341.845 7.77 341.975 ;
		RECT	14.68 341.845 14.73 341.975 ;
		RECT	9.1 339.195 9.15 339.325 ;
		RECT	10.81 339.195 10.86 339.325 ;
		RECT	9.1 341.615 9.15 341.745 ;
		RECT	10.81 341.615 10.86 341.745 ;
		RECT	6.76 342.075 6.81 342.205 ;
		RECT	8.04 342.075 8.09 342.205 ;
		RECT	9.58 342.075 9.63 342.205 ;
		RECT	9.855 342.075 9.905 342.205 ;
		RECT	10.26 342.075 10.31 342.205 ;
		RECT	11.565 342.075 11.615 342.205 ;
		RECT	13.33 342.075 13.38 342.205 ;
		RECT	6.765 344.495 6.815 344.625 ;
		RECT	8.04 344.495 8.09 344.625 ;
		RECT	9.58 344.495 9.63 344.625 ;
		RECT	9.855 344.495 9.905 344.625 ;
		RECT	11.565 344.495 11.615 344.625 ;
		RECT	13.33 344.495 13.38 344.625 ;
		RECT	7.72 344.725 7.77 344.855 ;
		RECT	14.68 344.725 14.73 344.855 ;
		RECT	9.1 342.075 9.15 342.205 ;
		RECT	10.81 342.075 10.86 342.205 ;
		RECT	9.1 344.495 9.15 344.625 ;
		RECT	10.81 344.495 10.86 344.625 ;
		RECT	6.76 344.955 6.81 345.085 ;
		RECT	8.04 344.955 8.09 345.085 ;
		RECT	9.58 344.955 9.63 345.085 ;
		RECT	9.855 344.955 9.905 345.085 ;
		RECT	10.26 344.955 10.31 345.085 ;
		RECT	11.565 344.955 11.615 345.085 ;
		RECT	13.33 344.955 13.38 345.085 ;
		RECT	6.765 347.375 6.815 347.505 ;
		RECT	8.04 347.375 8.09 347.505 ;
		RECT	9.58 347.375 9.63 347.505 ;
		RECT	9.855 347.375 9.905 347.505 ;
		RECT	11.565 347.375 11.615 347.505 ;
		RECT	13.33 347.375 13.38 347.505 ;
		RECT	7.72 347.605 7.77 347.735 ;
		RECT	14.68 347.605 14.73 347.735 ;
		RECT	9.1 344.955 9.15 345.085 ;
		RECT	10.81 344.955 10.86 345.085 ;
		RECT	9.1 347.375 9.15 347.505 ;
		RECT	10.81 347.375 10.86 347.505 ;
		RECT	6.76 347.835 6.81 347.965 ;
		RECT	8.04 347.835 8.09 347.965 ;
		RECT	9.58 347.835 9.63 347.965 ;
		RECT	9.855 347.835 9.905 347.965 ;
		RECT	10.26 347.835 10.31 347.965 ;
		RECT	11.565 347.835 11.615 347.965 ;
		RECT	13.33 347.835 13.38 347.965 ;
		RECT	6.765 350.255 6.815 350.385 ;
		RECT	8.04 350.255 8.09 350.385 ;
		RECT	9.58 350.255 9.63 350.385 ;
		RECT	9.855 350.255 9.905 350.385 ;
		RECT	11.565 350.255 11.615 350.385 ;
		RECT	13.33 350.255 13.38 350.385 ;
		RECT	7.72 350.485 7.77 350.615 ;
		RECT	14.68 350.485 14.73 350.615 ;
		RECT	9.1 347.835 9.15 347.965 ;
		RECT	10.81 347.835 10.86 347.965 ;
		RECT	9.1 350.255 9.15 350.385 ;
		RECT	10.81 350.255 10.86 350.385 ;
		RECT	6.76 350.715 6.81 350.845 ;
		RECT	8.04 350.715 8.09 350.845 ;
		RECT	9.58 350.715 9.63 350.845 ;
		RECT	9.855 350.715 9.905 350.845 ;
		RECT	10.26 350.715 10.31 350.845 ;
		RECT	11.565 350.715 11.615 350.845 ;
		RECT	13.33 350.715 13.38 350.845 ;
		RECT	6.765 353.135 6.815 353.265 ;
		RECT	8.04 353.135 8.09 353.265 ;
		RECT	9.58 353.135 9.63 353.265 ;
		RECT	9.855 353.135 9.905 353.265 ;
		RECT	11.565 353.135 11.615 353.265 ;
		RECT	13.33 353.135 13.38 353.265 ;
		RECT	7.72 353.365 7.77 353.495 ;
		RECT	14.68 353.365 14.73 353.495 ;
		RECT	9.1 350.715 9.15 350.845 ;
		RECT	10.81 350.715 10.86 350.845 ;
		RECT	9.1 353.135 9.15 353.265 ;
		RECT	10.81 353.135 10.86 353.265 ;
		RECT	6.76 353.595 6.81 353.725 ;
		RECT	8.04 353.595 8.09 353.725 ;
		RECT	9.58 353.595 9.63 353.725 ;
		RECT	9.855 353.595 9.905 353.725 ;
		RECT	10.26 353.595 10.31 353.725 ;
		RECT	11.565 353.595 11.615 353.725 ;
		RECT	13.33 353.595 13.38 353.725 ;
		RECT	6.765 356.015 6.815 356.145 ;
		RECT	8.04 356.015 8.09 356.145 ;
		RECT	9.58 356.015 9.63 356.145 ;
		RECT	9.855 356.015 9.905 356.145 ;
		RECT	11.565 356.015 11.615 356.145 ;
		RECT	13.33 356.015 13.38 356.145 ;
		RECT	7.72 356.245 7.77 356.375 ;
		RECT	14.68 356.245 14.73 356.375 ;
		RECT	9.1 353.595 9.15 353.725 ;
		RECT	10.81 353.595 10.86 353.725 ;
		RECT	9.1 356.015 9.15 356.145 ;
		RECT	10.81 356.015 10.86 356.145 ;
		RECT	6.76 356.475 6.81 356.605 ;
		RECT	8.04 356.475 8.09 356.605 ;
		RECT	9.58 356.475 9.63 356.605 ;
		RECT	9.855 356.475 9.905 356.605 ;
		RECT	10.26 356.475 10.31 356.605 ;
		RECT	11.565 356.475 11.615 356.605 ;
		RECT	13.33 356.475 13.38 356.605 ;
		RECT	6.765 358.895 6.815 359.025 ;
		RECT	8.04 358.895 8.09 359.025 ;
		RECT	9.58 358.895 9.63 359.025 ;
		RECT	9.855 358.895 9.905 359.025 ;
		RECT	11.565 358.895 11.615 359.025 ;
		RECT	13.33 358.895 13.38 359.025 ;
		RECT	7.72 359.125 7.77 359.255 ;
		RECT	14.68 359.125 14.73 359.255 ;
		RECT	9.1 356.475 9.15 356.605 ;
		RECT	10.81 356.475 10.86 356.605 ;
		RECT	9.1 358.895 9.15 359.025 ;
		RECT	10.81 358.895 10.86 359.025 ;
		RECT	6.76 359.355 6.81 359.485 ;
		RECT	8.04 359.355 8.09 359.485 ;
		RECT	9.58 359.355 9.63 359.485 ;
		RECT	9.855 359.355 9.905 359.485 ;
		RECT	10.26 359.355 10.31 359.485 ;
		RECT	11.565 359.355 11.615 359.485 ;
		RECT	13.33 359.355 13.38 359.485 ;
		RECT	6.765 361.775 6.815 361.905 ;
		RECT	8.04 361.775 8.09 361.905 ;
		RECT	9.58 361.775 9.63 361.905 ;
		RECT	9.855 361.775 9.905 361.905 ;
		RECT	11.565 361.775 11.615 361.905 ;
		RECT	13.33 361.775 13.38 361.905 ;
		RECT	7.72 362.005 7.77 362.135 ;
		RECT	14.68 362.005 14.73 362.135 ;
		RECT	9.1 359.355 9.15 359.485 ;
		RECT	10.81 359.355 10.86 359.485 ;
		RECT	9.1 361.775 9.15 361.905 ;
		RECT	10.81 361.775 10.86 361.905 ;
		RECT	6.76 362.235 6.81 362.365 ;
		RECT	8.04 362.235 8.09 362.365 ;
		RECT	9.58 362.235 9.63 362.365 ;
		RECT	9.855 362.235 9.905 362.365 ;
		RECT	10.26 362.235 10.31 362.365 ;
		RECT	11.565 362.235 11.615 362.365 ;
		RECT	13.33 362.235 13.38 362.365 ;
		RECT	6.765 364.655 6.815 364.785 ;
		RECT	8.04 364.655 8.09 364.785 ;
		RECT	9.58 364.655 9.63 364.785 ;
		RECT	9.855 364.655 9.905 364.785 ;
		RECT	11.565 364.655 11.615 364.785 ;
		RECT	13.33 364.655 13.38 364.785 ;
		RECT	7.72 364.885 7.77 365.015 ;
		RECT	14.68 364.885 14.73 365.015 ;
		RECT	9.1 362.235 9.15 362.365 ;
		RECT	10.81 362.235 10.86 362.365 ;
		RECT	9.1 364.655 9.15 364.785 ;
		RECT	10.81 364.655 10.86 364.785 ;
		RECT	6.76 365.115 6.81 365.245 ;
		RECT	8.04 365.115 8.09 365.245 ;
		RECT	9.58 365.115 9.63 365.245 ;
		RECT	9.855 365.115 9.905 365.245 ;
		RECT	10.26 365.115 10.31 365.245 ;
		RECT	11.565 365.115 11.615 365.245 ;
		RECT	13.33 365.115 13.38 365.245 ;
		RECT	6.765 367.535 6.815 367.665 ;
		RECT	8.04 367.535 8.09 367.665 ;
		RECT	9.58 367.535 9.63 367.665 ;
		RECT	9.855 367.535 9.905 367.665 ;
		RECT	11.565 367.535 11.615 367.665 ;
		RECT	13.33 367.535 13.38 367.665 ;
		RECT	7.72 367.765 7.77 367.895 ;
		RECT	14.68 367.765 14.73 367.895 ;
		RECT	9.1 365.115 9.15 365.245 ;
		RECT	10.81 365.115 10.86 365.245 ;
		RECT	9.1 367.535 9.15 367.665 ;
		RECT	10.81 367.535 10.86 367.665 ;
		RECT	6.76 367.995 6.81 368.125 ;
		RECT	8.04 367.995 8.09 368.125 ;
		RECT	9.58 367.995 9.63 368.125 ;
		RECT	9.855 367.995 9.905 368.125 ;
		RECT	10.26 367.995 10.31 368.125 ;
		RECT	11.565 367.995 11.615 368.125 ;
		RECT	13.33 367.995 13.38 368.125 ;
		RECT	6.765 370.415 6.815 370.545 ;
		RECT	8.04 370.415 8.09 370.545 ;
		RECT	9.58 370.415 9.63 370.545 ;
		RECT	9.855 370.415 9.905 370.545 ;
		RECT	11.565 370.415 11.615 370.545 ;
		RECT	13.33 370.415 13.38 370.545 ;
		RECT	7.72 370.645 7.77 370.775 ;
		RECT	14.68 370.645 14.73 370.775 ;
		RECT	9.1 367.995 9.15 368.125 ;
		RECT	10.81 367.995 10.86 368.125 ;
		RECT	9.1 370.415 9.15 370.545 ;
		RECT	10.81 370.415 10.86 370.545 ;
		RECT	6.76 370.875 6.81 371.005 ;
		RECT	8.04 370.875 8.09 371.005 ;
		RECT	9.58 370.875 9.63 371.005 ;
		RECT	9.855 370.875 9.905 371.005 ;
		RECT	10.26 370.875 10.31 371.005 ;
		RECT	11.565 370.875 11.615 371.005 ;
		RECT	13.33 370.875 13.38 371.005 ;
		RECT	6.765 373.295 6.815 373.425 ;
		RECT	8.04 373.295 8.09 373.425 ;
		RECT	9.58 373.295 9.63 373.425 ;
		RECT	9.855 373.295 9.905 373.425 ;
		RECT	11.565 373.295 11.615 373.425 ;
		RECT	13.33 373.295 13.38 373.425 ;
		RECT	7.72 373.525 7.77 373.655 ;
		RECT	14.68 373.525 14.73 373.655 ;
		RECT	9.1 370.875 9.15 371.005 ;
		RECT	10.81 370.875 10.86 371.005 ;
		RECT	9.1 373.295 9.15 373.425 ;
		RECT	10.81 373.295 10.86 373.425 ;
		RECT	6.76 373.755 6.81 373.885 ;
		RECT	8.04 373.755 8.09 373.885 ;
		RECT	9.58 373.755 9.63 373.885 ;
		RECT	9.855 373.755 9.905 373.885 ;
		RECT	10.26 373.755 10.31 373.885 ;
		RECT	11.565 373.755 11.615 373.885 ;
		RECT	13.33 373.755 13.38 373.885 ;
		RECT	6.765 376.175 6.815 376.305 ;
		RECT	8.04 376.175 8.09 376.305 ;
		RECT	9.58 376.175 9.63 376.305 ;
		RECT	9.855 376.175 9.905 376.305 ;
		RECT	11.565 376.175 11.615 376.305 ;
		RECT	13.33 376.175 13.38 376.305 ;
		RECT	7.72 376.405 7.77 376.535 ;
		RECT	14.68 376.405 14.73 376.535 ;
		RECT	9.1 373.755 9.15 373.885 ;
		RECT	10.81 373.755 10.86 373.885 ;
		RECT	9.1 376.175 9.15 376.305 ;
		RECT	10.81 376.175 10.86 376.305 ;
		RECT	6.76 376.635 6.81 376.765 ;
		RECT	8.04 376.635 8.09 376.765 ;
		RECT	9.58 376.635 9.63 376.765 ;
		RECT	9.855 376.635 9.905 376.765 ;
		RECT	10.26 376.635 10.31 376.765 ;
		RECT	11.565 376.635 11.615 376.765 ;
		RECT	13.33 376.635 13.38 376.765 ;
		RECT	6.765 379.055 6.815 379.185 ;
		RECT	8.04 379.055 8.09 379.185 ;
		RECT	9.58 379.055 9.63 379.185 ;
		RECT	9.855 379.055 9.905 379.185 ;
		RECT	11.565 379.055 11.615 379.185 ;
		RECT	13.33 379.055 13.38 379.185 ;
		RECT	7.72 379.285 7.77 379.415 ;
		RECT	14.68 379.285 14.73 379.415 ;
		RECT	9.1 376.635 9.15 376.765 ;
		RECT	10.81 376.635 10.86 376.765 ;
		RECT	9.1 379.055 9.15 379.185 ;
		RECT	10.81 379.055 10.86 379.185 ;
		RECT	6.76 379.515 6.81 379.645 ;
		RECT	8.04 379.515 8.09 379.645 ;
		RECT	9.58 379.515 9.63 379.645 ;
		RECT	9.855 379.515 9.905 379.645 ;
		RECT	10.26 379.515 10.31 379.645 ;
		RECT	11.565 379.515 11.615 379.645 ;
		RECT	13.33 379.515 13.38 379.645 ;
		RECT	6.765 381.935 6.815 382.065 ;
		RECT	8.04 381.935 8.09 382.065 ;
		RECT	9.58 381.935 9.63 382.065 ;
		RECT	9.855 381.935 9.905 382.065 ;
		RECT	11.565 381.935 11.615 382.065 ;
		RECT	13.33 381.935 13.38 382.065 ;
		RECT	7.72 382.165 7.77 382.295 ;
		RECT	14.68 382.165 14.73 382.295 ;
		RECT	9.1 379.515 9.15 379.645 ;
		RECT	10.81 379.515 10.86 379.645 ;
		RECT	9.1 381.935 9.15 382.065 ;
		RECT	10.81 381.935 10.86 382.065 ;
		RECT	6.76 382.395 6.81 382.525 ;
		RECT	8.04 382.395 8.09 382.525 ;
		RECT	9.58 382.395 9.63 382.525 ;
		RECT	9.855 382.395 9.905 382.525 ;
		RECT	10.26 382.395 10.31 382.525 ;
		RECT	11.565 382.395 11.615 382.525 ;
		RECT	13.33 382.395 13.38 382.525 ;
		RECT	6.765 384.815 6.815 384.945 ;
		RECT	8.04 384.815 8.09 384.945 ;
		RECT	9.58 384.815 9.63 384.945 ;
		RECT	9.855 384.815 9.905 384.945 ;
		RECT	11.565 384.815 11.615 384.945 ;
		RECT	13.33 384.815 13.38 384.945 ;
		RECT	7.72 385.045 7.77 385.175 ;
		RECT	14.68 385.045 14.73 385.175 ;
		RECT	9.1 382.395 9.15 382.525 ;
		RECT	10.81 382.395 10.86 382.525 ;
		RECT	9.1 384.815 9.15 384.945 ;
		RECT	10.81 384.815 10.86 384.945 ;
		RECT	6.76 385.275 6.81 385.405 ;
		RECT	8.04 385.275 8.09 385.405 ;
		RECT	9.58 385.275 9.63 385.405 ;
		RECT	9.855 385.275 9.905 385.405 ;
		RECT	10.26 385.275 10.31 385.405 ;
		RECT	11.565 385.275 11.615 385.405 ;
		RECT	13.33 385.275 13.38 385.405 ;
		RECT	6.765 387.695 6.815 387.825 ;
		RECT	8.04 387.695 8.09 387.825 ;
		RECT	9.58 387.695 9.63 387.825 ;
		RECT	9.855 387.695 9.905 387.825 ;
		RECT	11.565 387.695 11.615 387.825 ;
		RECT	13.33 387.695 13.38 387.825 ;
		RECT	7.72 387.925 7.77 388.055 ;
		RECT	14.68 387.925 14.73 388.055 ;
		RECT	9.1 385.275 9.15 385.405 ;
		RECT	10.81 385.275 10.86 385.405 ;
		RECT	9.1 387.695 9.15 387.825 ;
		RECT	10.81 387.695 10.86 387.825 ;
		RECT	6.76 388.155 6.81 388.285 ;
		RECT	8.04 388.155 8.09 388.285 ;
		RECT	9.58 388.155 9.63 388.285 ;
		RECT	9.855 388.155 9.905 388.285 ;
		RECT	10.26 388.155 10.31 388.285 ;
		RECT	11.565 388.155 11.615 388.285 ;
		RECT	13.33 388.155 13.38 388.285 ;
		RECT	6.765 390.575 6.815 390.705 ;
		RECT	8.04 390.575 8.09 390.705 ;
		RECT	9.58 390.575 9.63 390.705 ;
		RECT	9.855 390.575 9.905 390.705 ;
		RECT	11.565 390.575 11.615 390.705 ;
		RECT	13.33 390.575 13.38 390.705 ;
		RECT	7.72 390.805 7.77 390.935 ;
		RECT	14.68 390.805 14.73 390.935 ;
		RECT	9.1 388.155 9.15 388.285 ;
		RECT	10.81 388.155 10.86 388.285 ;
		RECT	9.1 390.575 9.15 390.705 ;
		RECT	10.81 390.575 10.86 390.705 ;
		RECT	6.76 391.035 6.81 391.165 ;
		RECT	8.04 391.035 8.09 391.165 ;
		RECT	9.58 391.035 9.63 391.165 ;
		RECT	9.855 391.035 9.905 391.165 ;
		RECT	10.26 391.035 10.31 391.165 ;
		RECT	11.565 391.035 11.615 391.165 ;
		RECT	13.33 391.035 13.38 391.165 ;
		RECT	6.765 393.455 6.815 393.585 ;
		RECT	8.04 393.455 8.09 393.585 ;
		RECT	9.58 393.455 9.63 393.585 ;
		RECT	9.855 393.455 9.905 393.585 ;
		RECT	11.565 393.455 11.615 393.585 ;
		RECT	13.33 393.455 13.38 393.585 ;
		RECT	7.72 393.685 7.77 393.815 ;
		RECT	14.68 393.685 14.73 393.815 ;
		RECT	9.1 391.035 9.15 391.165 ;
		RECT	10.81 391.035 10.86 391.165 ;
		RECT	9.1 393.455 9.15 393.585 ;
		RECT	10.81 393.455 10.86 393.585 ;
		RECT	6.76 393.915 6.81 394.045 ;
		RECT	8.04 393.915 8.09 394.045 ;
		RECT	9.58 393.915 9.63 394.045 ;
		RECT	9.855 393.915 9.905 394.045 ;
		RECT	10.26 393.915 10.31 394.045 ;
		RECT	11.565 393.915 11.615 394.045 ;
		RECT	13.33 393.915 13.38 394.045 ;
		RECT	6.765 396.335 6.815 396.465 ;
		RECT	8.04 396.335 8.09 396.465 ;
		RECT	9.58 396.335 9.63 396.465 ;
		RECT	9.855 396.335 9.905 396.465 ;
		RECT	11.565 396.335 11.615 396.465 ;
		RECT	13.33 396.335 13.38 396.465 ;
		RECT	7.72 396.565 7.77 396.695 ;
		RECT	14.68 396.565 14.73 396.695 ;
		RECT	9.1 393.915 9.15 394.045 ;
		RECT	10.81 393.915 10.86 394.045 ;
		RECT	9.1 396.335 9.15 396.465 ;
		RECT	10.81 396.335 10.86 396.465 ;
		RECT	6.76 396.795 6.81 396.925 ;
		RECT	8.04 396.795 8.09 396.925 ;
		RECT	9.58 396.795 9.63 396.925 ;
		RECT	9.855 396.795 9.905 396.925 ;
		RECT	10.26 396.795 10.31 396.925 ;
		RECT	11.565 396.795 11.615 396.925 ;
		RECT	13.33 396.795 13.38 396.925 ;
		RECT	6.765 399.215 6.815 399.345 ;
		RECT	8.04 399.215 8.09 399.345 ;
		RECT	9.58 399.215 9.63 399.345 ;
		RECT	9.855 399.215 9.905 399.345 ;
		RECT	11.565 399.215 11.615 399.345 ;
		RECT	13.33 399.215 13.38 399.345 ;
		RECT	7.72 399.445 7.77 399.575 ;
		RECT	14.68 399.445 14.73 399.575 ;
		RECT	9.1 396.795 9.15 396.925 ;
		RECT	10.81 396.795 10.86 396.925 ;
		RECT	9.1 399.215 9.15 399.345 ;
		RECT	10.81 399.215 10.86 399.345 ;
		RECT	6.76 399.675 6.81 399.805 ;
		RECT	8.04 399.675 8.09 399.805 ;
		RECT	9.58 399.675 9.63 399.805 ;
		RECT	9.855 399.675 9.905 399.805 ;
		RECT	10.26 399.675 10.31 399.805 ;
		RECT	11.565 399.675 11.615 399.805 ;
		RECT	13.33 399.675 13.38 399.805 ;
		RECT	6.765 402.095 6.815 402.225 ;
		RECT	8.04 402.095 8.09 402.225 ;
		RECT	9.58 402.095 9.63 402.225 ;
		RECT	9.855 402.095 9.905 402.225 ;
		RECT	11.565 402.095 11.615 402.225 ;
		RECT	13.33 402.095 13.38 402.225 ;
		RECT	7.72 402.325 7.77 402.455 ;
		RECT	14.68 402.325 14.73 402.455 ;
		RECT	9.1 399.675 9.15 399.805 ;
		RECT	10.81 399.675 10.86 399.805 ;
		RECT	9.1 402.095 9.15 402.225 ;
		RECT	10.81 402.095 10.86 402.225 ;
		RECT	6.76 402.555 6.81 402.685 ;
		RECT	8.04 402.555 8.09 402.685 ;
		RECT	9.58 402.555 9.63 402.685 ;
		RECT	9.855 402.555 9.905 402.685 ;
		RECT	10.26 402.555 10.31 402.685 ;
		RECT	11.565 402.555 11.615 402.685 ;
		RECT	13.33 402.555 13.38 402.685 ;
		RECT	6.765 404.975 6.815 405.105 ;
		RECT	8.04 404.975 8.09 405.105 ;
		RECT	9.58 404.975 9.63 405.105 ;
		RECT	9.855 404.975 9.905 405.105 ;
		RECT	11.565 404.975 11.615 405.105 ;
		RECT	13.33 404.975 13.38 405.105 ;
		RECT	7.72 405.205 7.77 405.335 ;
		RECT	14.68 405.205 14.73 405.335 ;
		RECT	9.1 402.555 9.15 402.685 ;
		RECT	10.81 402.555 10.86 402.685 ;
		RECT	9.1 404.975 9.15 405.105 ;
		RECT	10.81 404.975 10.86 405.105 ;
		RECT	6.76 405.435 6.81 405.565 ;
		RECT	8.04 405.435 8.09 405.565 ;
		RECT	9.58 405.435 9.63 405.565 ;
		RECT	9.855 405.435 9.905 405.565 ;
		RECT	10.26 405.435 10.31 405.565 ;
		RECT	11.565 405.435 11.615 405.565 ;
		RECT	13.33 405.435 13.38 405.565 ;
		RECT	6.765 407.855 6.815 407.985 ;
		RECT	8.04 407.855 8.09 407.985 ;
		RECT	9.58 407.855 9.63 407.985 ;
		RECT	9.855 407.855 9.905 407.985 ;
		RECT	11.565 407.855 11.615 407.985 ;
		RECT	13.33 407.855 13.38 407.985 ;
		RECT	7.72 408.085 7.77 408.215 ;
		RECT	14.68 408.085 14.73 408.215 ;
		RECT	9.1 405.435 9.15 405.565 ;
		RECT	10.81 405.435 10.86 405.565 ;
		RECT	9.1 407.855 9.15 407.985 ;
		RECT	10.81 407.855 10.86 407.985 ;
		RECT	6.76 408.315 6.81 408.445 ;
		RECT	8.04 408.315 8.09 408.445 ;
		RECT	9.58 408.315 9.63 408.445 ;
		RECT	9.855 408.315 9.905 408.445 ;
		RECT	10.26 408.315 10.31 408.445 ;
		RECT	11.565 408.315 11.615 408.445 ;
		RECT	13.33 408.315 13.38 408.445 ;
		RECT	6.765 410.735 6.815 410.865 ;
		RECT	8.04 410.735 8.09 410.865 ;
		RECT	9.58 410.735 9.63 410.865 ;
		RECT	9.855 410.735 9.905 410.865 ;
		RECT	11.565 410.735 11.615 410.865 ;
		RECT	13.33 410.735 13.38 410.865 ;
		RECT	7.72 410.965 7.77 411.095 ;
		RECT	14.68 410.965 14.73 411.095 ;
		RECT	9.1 408.315 9.15 408.445 ;
		RECT	10.81 408.315 10.86 408.445 ;
		RECT	9.1 410.735 9.15 410.865 ;
		RECT	10.81 410.735 10.86 410.865 ;
		RECT	6.76 411.195 6.81 411.325 ;
		RECT	8.04 411.195 8.09 411.325 ;
		RECT	9.58 411.195 9.63 411.325 ;
		RECT	9.855 411.195 9.905 411.325 ;
		RECT	10.26 411.195 10.31 411.325 ;
		RECT	11.565 411.195 11.615 411.325 ;
		RECT	13.33 411.195 13.38 411.325 ;
		RECT	6.765 413.615 6.815 413.745 ;
		RECT	8.04 413.615 8.09 413.745 ;
		RECT	9.58 413.615 9.63 413.745 ;
		RECT	9.855 413.615 9.905 413.745 ;
		RECT	11.565 413.615 11.615 413.745 ;
		RECT	13.33 413.615 13.38 413.745 ;
		RECT	7.72 413.845 7.77 413.975 ;
		RECT	14.68 413.845 14.73 413.975 ;
		RECT	9.1 411.195 9.15 411.325 ;
		RECT	10.81 411.195 10.86 411.325 ;
		RECT	9.1 413.615 9.15 413.745 ;
		RECT	10.81 413.615 10.86 413.745 ;
		RECT	14.87 232.635 14.92 232.765 ;
		RECT	6.76 233.095 6.81 233.225 ;
		RECT	8.04 233.095 8.09 233.225 ;
		RECT	9.58 233.095 9.63 233.225 ;
		RECT	9.855 233.095 9.905 233.225 ;
		RECT	10.26 233.095 10.31 233.225 ;
		RECT	11.565 233.095 11.615 233.225 ;
		RECT	13.33 233.095 13.38 233.225 ;
		RECT	14.23 233.095 14.28 233.225 ;
		RECT	14.23 234.825 14.28 234.955 ;
		RECT	14.87 235.055 14.92 235.185 ;
		RECT	6.215 235.285 6.265 235.415 ;
		RECT	6.605 235.285 6.655 235.415 ;
		RECT	7.265 235.285 7.315 235.415 ;
		RECT	8.96 235.285 9.01 235.415 ;
		RECT	9.31 235.285 9.36 235.415 ;
		RECT	12.095 235.285 12.145 235.415 ;
		RECT	12.355 235.285 12.405 235.415 ;
		RECT	13.06 235.285 13.11 235.415 ;
		RECT	14.52 235.285 14.57 235.415 ;
		RECT	14.87 258.555 14.92 258.685 ;
		RECT	6.76 259.015 6.81 259.145 ;
		RECT	8.04 259.015 8.09 259.145 ;
		RECT	9.58 259.015 9.63 259.145 ;
		RECT	9.855 259.015 9.905 259.145 ;
		RECT	10.26 259.015 10.31 259.145 ;
		RECT	11.565 259.015 11.615 259.145 ;
		RECT	13.33 259.015 13.38 259.145 ;
		RECT	14.23 259.015 14.28 259.145 ;
		RECT	14.23 260.745 14.28 260.875 ;
		RECT	14.87 260.975 14.92 261.105 ;
		RECT	6.215 261.205 6.265 261.335 ;
		RECT	6.605 261.205 6.655 261.335 ;
		RECT	7.265 261.205 7.315 261.335 ;
		RECT	8.96 261.205 9.01 261.335 ;
		RECT	9.31 261.205 9.36 261.335 ;
		RECT	12.095 261.205 12.145 261.335 ;
		RECT	12.355 261.205 12.405 261.335 ;
		RECT	13.06 261.205 13.11 261.335 ;
		RECT	14.52 261.205 14.57 261.335 ;
		RECT	14.87 261.435 14.92 261.565 ;
		RECT	6.76 261.895 6.81 262.025 ;
		RECT	8.04 261.895 8.09 262.025 ;
		RECT	9.58 261.895 9.63 262.025 ;
		RECT	9.855 261.895 9.905 262.025 ;
		RECT	10.26 261.895 10.31 262.025 ;
		RECT	11.565 261.895 11.615 262.025 ;
		RECT	13.33 261.895 13.38 262.025 ;
		RECT	14.23 261.895 14.28 262.025 ;
		RECT	14.23 263.625 14.28 263.755 ;
		RECT	14.87 263.855 14.92 263.985 ;
		RECT	6.215 264.085 6.265 264.215 ;
		RECT	6.605 264.085 6.655 264.215 ;
		RECT	7.265 264.085 7.315 264.215 ;
		RECT	8.96 264.085 9.01 264.215 ;
		RECT	9.31 264.085 9.36 264.215 ;
		RECT	12.095 264.085 12.145 264.215 ;
		RECT	12.355 264.085 12.405 264.215 ;
		RECT	13.06 264.085 13.11 264.215 ;
		RECT	14.52 264.085 14.57 264.215 ;
		RECT	14.87 264.315 14.92 264.445 ;
		RECT	6.76 264.775 6.81 264.905 ;
		RECT	8.04 264.775 8.09 264.905 ;
		RECT	9.58 264.775 9.63 264.905 ;
		RECT	9.855 264.775 9.905 264.905 ;
		RECT	10.26 264.775 10.31 264.905 ;
		RECT	11.565 264.775 11.615 264.905 ;
		RECT	13.33 264.775 13.38 264.905 ;
		RECT	14.23 264.775 14.28 264.905 ;
		RECT	14.23 266.505 14.28 266.635 ;
		RECT	14.87 266.735 14.92 266.865 ;
		RECT	6.215 266.965 6.265 267.095 ;
		RECT	6.605 266.965 6.655 267.095 ;
		RECT	7.265 266.965 7.315 267.095 ;
		RECT	8.96 266.965 9.01 267.095 ;
		RECT	9.31 266.965 9.36 267.095 ;
		RECT	12.095 266.965 12.145 267.095 ;
		RECT	12.355 266.965 12.405 267.095 ;
		RECT	13.06 266.965 13.11 267.095 ;
		RECT	14.52 266.965 14.57 267.095 ;
		RECT	14.87 267.195 14.92 267.325 ;
		RECT	6.76 267.655 6.81 267.785 ;
		RECT	8.04 267.655 8.09 267.785 ;
		RECT	9.58 267.655 9.63 267.785 ;
		RECT	9.855 267.655 9.905 267.785 ;
		RECT	10.26 267.655 10.31 267.785 ;
		RECT	11.565 267.655 11.615 267.785 ;
		RECT	13.33 267.655 13.38 267.785 ;
		RECT	14.23 267.655 14.28 267.785 ;
		RECT	14.23 269.385 14.28 269.515 ;
		RECT	14.87 269.615 14.92 269.745 ;
		RECT	6.215 269.845 6.265 269.975 ;
		RECT	6.605 269.845 6.655 269.975 ;
		RECT	7.265 269.845 7.315 269.975 ;
		RECT	8.96 269.845 9.01 269.975 ;
		RECT	9.31 269.845 9.36 269.975 ;
		RECT	12.095 269.845 12.145 269.975 ;
		RECT	12.355 269.845 12.405 269.975 ;
		RECT	13.06 269.845 13.11 269.975 ;
		RECT	14.52 269.845 14.57 269.975 ;
		RECT	14.87 270.075 14.92 270.205 ;
		RECT	6.76 270.535 6.81 270.665 ;
		RECT	8.04 270.535 8.09 270.665 ;
		RECT	9.58 270.535 9.63 270.665 ;
		RECT	9.855 270.535 9.905 270.665 ;
		RECT	10.26 270.535 10.31 270.665 ;
		RECT	11.565 270.535 11.615 270.665 ;
		RECT	13.33 270.535 13.38 270.665 ;
		RECT	14.23 270.535 14.28 270.665 ;
		RECT	14.23 272.265 14.28 272.395 ;
		RECT	14.87 272.495 14.92 272.625 ;
		RECT	6.215 272.725 6.265 272.855 ;
		RECT	6.605 272.725 6.655 272.855 ;
		RECT	7.265 272.725 7.315 272.855 ;
		RECT	8.96 272.725 9.01 272.855 ;
		RECT	9.31 272.725 9.36 272.855 ;
		RECT	12.095 272.725 12.145 272.855 ;
		RECT	12.355 272.725 12.405 272.855 ;
		RECT	13.06 272.725 13.11 272.855 ;
		RECT	14.52 272.725 14.57 272.855 ;
		RECT	14.87 272.955 14.92 273.085 ;
		RECT	6.76 273.415 6.81 273.545 ;
		RECT	8.04 273.415 8.09 273.545 ;
		RECT	9.58 273.415 9.63 273.545 ;
		RECT	9.855 273.415 9.905 273.545 ;
		RECT	10.26 273.415 10.31 273.545 ;
		RECT	11.565 273.415 11.615 273.545 ;
		RECT	13.33 273.415 13.38 273.545 ;
		RECT	14.23 273.415 14.28 273.545 ;
		RECT	14.23 275.145 14.28 275.275 ;
		RECT	14.87 275.375 14.92 275.505 ;
		RECT	6.215 275.605 6.265 275.735 ;
		RECT	6.605 275.605 6.655 275.735 ;
		RECT	7.265 275.605 7.315 275.735 ;
		RECT	8.96 275.605 9.01 275.735 ;
		RECT	9.31 275.605 9.36 275.735 ;
		RECT	12.095 275.605 12.145 275.735 ;
		RECT	12.355 275.605 12.405 275.735 ;
		RECT	13.06 275.605 13.11 275.735 ;
		RECT	14.52 275.605 14.57 275.735 ;
		RECT	14.87 275.835 14.92 275.965 ;
		RECT	6.76 276.295 6.81 276.425 ;
		RECT	8.04 276.295 8.09 276.425 ;
		RECT	9.58 276.295 9.63 276.425 ;
		RECT	9.855 276.295 9.905 276.425 ;
		RECT	10.26 276.295 10.31 276.425 ;
		RECT	11.565 276.295 11.615 276.425 ;
		RECT	13.33 276.295 13.38 276.425 ;
		RECT	14.23 276.295 14.28 276.425 ;
		RECT	14.23 278.025 14.28 278.155 ;
		RECT	14.87 278.255 14.92 278.385 ;
		RECT	6.215 278.485 6.265 278.615 ;
		RECT	6.605 278.485 6.655 278.615 ;
		RECT	7.265 278.485 7.315 278.615 ;
		RECT	8.96 278.485 9.01 278.615 ;
		RECT	9.31 278.485 9.36 278.615 ;
		RECT	12.095 278.485 12.145 278.615 ;
		RECT	12.355 278.485 12.405 278.615 ;
		RECT	13.06 278.485 13.11 278.615 ;
		RECT	14.52 278.485 14.57 278.615 ;
		RECT	14.87 278.715 14.92 278.845 ;
		RECT	6.76 279.175 6.81 279.305 ;
		RECT	8.04 279.175 8.09 279.305 ;
		RECT	9.58 279.175 9.63 279.305 ;
		RECT	9.855 279.175 9.905 279.305 ;
		RECT	10.26 279.175 10.31 279.305 ;
		RECT	11.565 279.175 11.615 279.305 ;
		RECT	13.33 279.175 13.38 279.305 ;
		RECT	14.23 279.175 14.28 279.305 ;
		RECT	14.23 280.905 14.28 281.035 ;
		RECT	14.87 281.135 14.92 281.265 ;
		RECT	6.215 281.365 6.265 281.495 ;
		RECT	6.605 281.365 6.655 281.495 ;
		RECT	7.265 281.365 7.315 281.495 ;
		RECT	8.96 281.365 9.01 281.495 ;
		RECT	9.31 281.365 9.36 281.495 ;
		RECT	12.095 281.365 12.145 281.495 ;
		RECT	12.355 281.365 12.405 281.495 ;
		RECT	13.06 281.365 13.11 281.495 ;
		RECT	14.52 281.365 14.57 281.495 ;
		RECT	14.87 281.595 14.92 281.725 ;
		RECT	6.76 282.055 6.81 282.185 ;
		RECT	8.04 282.055 8.09 282.185 ;
		RECT	9.58 282.055 9.63 282.185 ;
		RECT	9.855 282.055 9.905 282.185 ;
		RECT	10.26 282.055 10.31 282.185 ;
		RECT	11.565 282.055 11.615 282.185 ;
		RECT	13.33 282.055 13.38 282.185 ;
		RECT	14.23 282.055 14.28 282.185 ;
		RECT	14.23 283.785 14.28 283.915 ;
		RECT	14.87 284.015 14.92 284.145 ;
		RECT	6.215 284.245 6.265 284.375 ;
		RECT	6.605 284.245 6.655 284.375 ;
		RECT	7.265 284.245 7.315 284.375 ;
		RECT	8.96 284.245 9.01 284.375 ;
		RECT	9.31 284.245 9.36 284.375 ;
		RECT	12.095 284.245 12.145 284.375 ;
		RECT	12.355 284.245 12.405 284.375 ;
		RECT	13.06 284.245 13.11 284.375 ;
		RECT	14.52 284.245 14.57 284.375 ;
		RECT	14.87 284.475 14.92 284.605 ;
		RECT	6.76 284.935 6.81 285.065 ;
		RECT	8.04 284.935 8.09 285.065 ;
		RECT	9.58 284.935 9.63 285.065 ;
		RECT	9.855 284.935 9.905 285.065 ;
		RECT	10.26 284.935 10.31 285.065 ;
		RECT	11.565 284.935 11.615 285.065 ;
		RECT	13.33 284.935 13.38 285.065 ;
		RECT	14.23 284.935 14.28 285.065 ;
		RECT	14.23 286.665 14.28 286.795 ;
		RECT	14.87 286.895 14.92 287.025 ;
		RECT	6.215 287.125 6.265 287.255 ;
		RECT	6.605 287.125 6.655 287.255 ;
		RECT	7.265 287.125 7.315 287.255 ;
		RECT	8.96 287.125 9.01 287.255 ;
		RECT	9.31 287.125 9.36 287.255 ;
		RECT	12.095 287.125 12.145 287.255 ;
		RECT	12.355 287.125 12.405 287.255 ;
		RECT	13.06 287.125 13.11 287.255 ;
		RECT	14.52 287.125 14.57 287.255 ;
		RECT	14.87 235.515 14.92 235.645 ;
		RECT	6.76 235.975 6.81 236.105 ;
		RECT	8.04 235.975 8.09 236.105 ;
		RECT	9.58 235.975 9.63 236.105 ;
		RECT	9.855 235.975 9.905 236.105 ;
		RECT	10.26 235.975 10.31 236.105 ;
		RECT	11.565 235.975 11.615 236.105 ;
		RECT	13.33 235.975 13.38 236.105 ;
		RECT	14.23 235.975 14.28 236.105 ;
		RECT	14.23 237.705 14.28 237.835 ;
		RECT	14.87 237.935 14.92 238.065 ;
		RECT	6.215 238.165 6.265 238.295 ;
		RECT	6.605 238.165 6.655 238.295 ;
		RECT	7.265 238.165 7.315 238.295 ;
		RECT	8.96 238.165 9.01 238.295 ;
		RECT	9.31 238.165 9.36 238.295 ;
		RECT	12.095 238.165 12.145 238.295 ;
		RECT	12.355 238.165 12.405 238.295 ;
		RECT	13.06 238.165 13.11 238.295 ;
		RECT	14.52 238.165 14.57 238.295 ;
		RECT	14.87 287.355 14.92 287.485 ;
		RECT	6.76 287.815 6.81 287.945 ;
		RECT	8.04 287.815 8.09 287.945 ;
		RECT	9.58 287.815 9.63 287.945 ;
		RECT	9.855 287.815 9.905 287.945 ;
		RECT	10.26 287.815 10.31 287.945 ;
		RECT	11.565 287.815 11.615 287.945 ;
		RECT	13.33 287.815 13.38 287.945 ;
		RECT	14.23 287.815 14.28 287.945 ;
		RECT	14.23 289.545 14.28 289.675 ;
		RECT	14.87 289.775 14.92 289.905 ;
		RECT	6.215 290.005 6.265 290.135 ;
		RECT	6.605 290.005 6.655 290.135 ;
		RECT	7.265 290.005 7.315 290.135 ;
		RECT	8.96 290.005 9.01 290.135 ;
		RECT	9.31 290.005 9.36 290.135 ;
		RECT	12.095 290.005 12.145 290.135 ;
		RECT	12.355 290.005 12.405 290.135 ;
		RECT	13.06 290.005 13.11 290.135 ;
		RECT	14.52 290.005 14.57 290.135 ;
		RECT	14.87 290.235 14.92 290.365 ;
		RECT	6.76 290.695 6.81 290.825 ;
		RECT	8.04 290.695 8.09 290.825 ;
		RECT	9.58 290.695 9.63 290.825 ;
		RECT	9.855 290.695 9.905 290.825 ;
		RECT	10.26 290.695 10.31 290.825 ;
		RECT	11.565 290.695 11.615 290.825 ;
		RECT	13.33 290.695 13.38 290.825 ;
		RECT	14.23 290.695 14.28 290.825 ;
		RECT	14.23 292.425 14.28 292.555 ;
		RECT	14.87 292.655 14.92 292.785 ;
		RECT	6.215 292.885 6.265 293.015 ;
		RECT	6.605 292.885 6.655 293.015 ;
		RECT	7.265 292.885 7.315 293.015 ;
		RECT	8.96 292.885 9.01 293.015 ;
		RECT	9.31 292.885 9.36 293.015 ;
		RECT	12.095 292.885 12.145 293.015 ;
		RECT	12.355 292.885 12.405 293.015 ;
		RECT	13.06 292.885 13.11 293.015 ;
		RECT	14.52 292.885 14.57 293.015 ;
		RECT	14.87 293.115 14.92 293.245 ;
		RECT	6.76 293.575 6.81 293.705 ;
		RECT	8.04 293.575 8.09 293.705 ;
		RECT	9.58 293.575 9.63 293.705 ;
		RECT	9.855 293.575 9.905 293.705 ;
		RECT	10.26 293.575 10.31 293.705 ;
		RECT	11.565 293.575 11.615 293.705 ;
		RECT	13.33 293.575 13.38 293.705 ;
		RECT	14.23 293.575 14.28 293.705 ;
		RECT	14.23 295.305 14.28 295.435 ;
		RECT	14.87 295.535 14.92 295.665 ;
		RECT	6.215 295.765 6.265 295.895 ;
		RECT	6.605 295.765 6.655 295.895 ;
		RECT	7.265 295.765 7.315 295.895 ;
		RECT	8.96 295.765 9.01 295.895 ;
		RECT	9.31 295.765 9.36 295.895 ;
		RECT	12.095 295.765 12.145 295.895 ;
		RECT	12.355 295.765 12.405 295.895 ;
		RECT	13.06 295.765 13.11 295.895 ;
		RECT	14.52 295.765 14.57 295.895 ;
		RECT	14.87 295.995 14.92 296.125 ;
		RECT	6.76 296.455 6.81 296.585 ;
		RECT	8.04 296.455 8.09 296.585 ;
		RECT	9.58 296.455 9.63 296.585 ;
		RECT	9.855 296.455 9.905 296.585 ;
		RECT	10.26 296.455 10.31 296.585 ;
		RECT	11.565 296.455 11.615 296.585 ;
		RECT	13.33 296.455 13.38 296.585 ;
		RECT	14.23 296.455 14.28 296.585 ;
		RECT	14.23 298.185 14.28 298.315 ;
		RECT	14.87 298.415 14.92 298.545 ;
		RECT	6.215 298.645 6.265 298.775 ;
		RECT	6.605 298.645 6.655 298.775 ;
		RECT	7.265 298.645 7.315 298.775 ;
		RECT	8.96 298.645 9.01 298.775 ;
		RECT	9.31 298.645 9.36 298.775 ;
		RECT	12.095 298.645 12.145 298.775 ;
		RECT	12.355 298.645 12.405 298.775 ;
		RECT	13.06 298.645 13.11 298.775 ;
		RECT	14.52 298.645 14.57 298.775 ;
		RECT	14.87 298.875 14.92 299.005 ;
		RECT	6.76 299.335 6.81 299.465 ;
		RECT	8.04 299.335 8.09 299.465 ;
		RECT	9.58 299.335 9.63 299.465 ;
		RECT	9.855 299.335 9.905 299.465 ;
		RECT	10.26 299.335 10.31 299.465 ;
		RECT	11.565 299.335 11.615 299.465 ;
		RECT	13.33 299.335 13.38 299.465 ;
		RECT	14.23 299.335 14.28 299.465 ;
		RECT	14.23 301.065 14.28 301.195 ;
		RECT	14.87 301.295 14.92 301.425 ;
		RECT	6.215 301.525 6.265 301.655 ;
		RECT	6.605 301.525 6.655 301.655 ;
		RECT	7.265 301.525 7.315 301.655 ;
		RECT	8.96 301.525 9.01 301.655 ;
		RECT	9.31 301.525 9.36 301.655 ;
		RECT	12.095 301.525 12.145 301.655 ;
		RECT	12.355 301.525 12.405 301.655 ;
		RECT	13.06 301.525 13.11 301.655 ;
		RECT	14.52 301.525 14.57 301.655 ;
		RECT	14.87 301.755 14.92 301.885 ;
		RECT	6.76 302.215 6.81 302.345 ;
		RECT	8.04 302.215 8.09 302.345 ;
		RECT	9.58 302.215 9.63 302.345 ;
		RECT	9.855 302.215 9.905 302.345 ;
		RECT	10.26 302.215 10.31 302.345 ;
		RECT	11.565 302.215 11.615 302.345 ;
		RECT	13.33 302.215 13.38 302.345 ;
		RECT	14.23 302.215 14.28 302.345 ;
		RECT	14.23 303.945 14.28 304.075 ;
		RECT	14.87 304.175 14.92 304.305 ;
		RECT	6.215 304.405 6.265 304.535 ;
		RECT	6.605 304.405 6.655 304.535 ;
		RECT	7.265 304.405 7.315 304.535 ;
		RECT	8.96 304.405 9.01 304.535 ;
		RECT	9.31 304.405 9.36 304.535 ;
		RECT	12.095 304.405 12.145 304.535 ;
		RECT	12.355 304.405 12.405 304.535 ;
		RECT	13.06 304.405 13.11 304.535 ;
		RECT	14.52 304.405 14.57 304.535 ;
		RECT	14.87 304.635 14.92 304.765 ;
		RECT	6.76 305.095 6.81 305.225 ;
		RECT	8.04 305.095 8.09 305.225 ;
		RECT	9.58 305.095 9.63 305.225 ;
		RECT	9.855 305.095 9.905 305.225 ;
		RECT	10.26 305.095 10.31 305.225 ;
		RECT	11.565 305.095 11.615 305.225 ;
		RECT	13.33 305.095 13.38 305.225 ;
		RECT	14.23 305.095 14.28 305.225 ;
		RECT	14.23 306.825 14.28 306.955 ;
		RECT	14.87 307.055 14.92 307.185 ;
		RECT	6.215 307.285 6.265 307.415 ;
		RECT	6.605 307.285 6.655 307.415 ;
		RECT	7.265 307.285 7.315 307.415 ;
		RECT	8.96 307.285 9.01 307.415 ;
		RECT	9.31 307.285 9.36 307.415 ;
		RECT	12.095 307.285 12.145 307.415 ;
		RECT	12.355 307.285 12.405 307.415 ;
		RECT	13.06 307.285 13.11 307.415 ;
		RECT	14.52 307.285 14.57 307.415 ;
		RECT	14.87 307.515 14.92 307.645 ;
		RECT	6.76 307.975 6.81 308.105 ;
		RECT	8.04 307.975 8.09 308.105 ;
		RECT	9.58 307.975 9.63 308.105 ;
		RECT	9.855 307.975 9.905 308.105 ;
		RECT	10.26 307.975 10.31 308.105 ;
		RECT	11.565 307.975 11.615 308.105 ;
		RECT	13.33 307.975 13.38 308.105 ;
		RECT	14.23 307.975 14.28 308.105 ;
		RECT	14.23 309.705 14.28 309.835 ;
		RECT	14.87 309.935 14.92 310.065 ;
		RECT	6.215 310.165 6.265 310.295 ;
		RECT	6.605 310.165 6.655 310.295 ;
		RECT	7.265 310.165 7.315 310.295 ;
		RECT	8.96 310.165 9.01 310.295 ;
		RECT	9.31 310.165 9.36 310.295 ;
		RECT	12.095 310.165 12.145 310.295 ;
		RECT	12.355 310.165 12.405 310.295 ;
		RECT	13.06 310.165 13.11 310.295 ;
		RECT	14.52 310.165 14.57 310.295 ;
		RECT	14.87 310.395 14.92 310.525 ;
		RECT	6.76 310.855 6.81 310.985 ;
		RECT	8.04 310.855 8.09 310.985 ;
		RECT	9.58 310.855 9.63 310.985 ;
		RECT	9.855 310.855 9.905 310.985 ;
		RECT	10.26 310.855 10.31 310.985 ;
		RECT	11.565 310.855 11.615 310.985 ;
		RECT	13.33 310.855 13.38 310.985 ;
		RECT	14.23 310.855 14.28 310.985 ;
		RECT	14.23 312.585 14.28 312.715 ;
		RECT	14.87 312.815 14.92 312.945 ;
		RECT	6.215 313.045 6.265 313.175 ;
		RECT	6.605 313.045 6.655 313.175 ;
		RECT	7.265 313.045 7.315 313.175 ;
		RECT	8.96 313.045 9.01 313.175 ;
		RECT	9.31 313.045 9.36 313.175 ;
		RECT	12.095 313.045 12.145 313.175 ;
		RECT	12.355 313.045 12.405 313.175 ;
		RECT	13.06 313.045 13.11 313.175 ;
		RECT	14.52 313.045 14.57 313.175 ;
		RECT	14.87 313.275 14.92 313.405 ;
		RECT	6.76 313.735 6.81 313.865 ;
		RECT	8.04 313.735 8.09 313.865 ;
		RECT	9.58 313.735 9.63 313.865 ;
		RECT	9.855 313.735 9.905 313.865 ;
		RECT	10.26 313.735 10.31 313.865 ;
		RECT	11.565 313.735 11.615 313.865 ;
		RECT	13.33 313.735 13.38 313.865 ;
		RECT	14.23 313.735 14.28 313.865 ;
		RECT	14.23 315.465 14.28 315.595 ;
		RECT	14.87 315.695 14.92 315.825 ;
		RECT	6.215 315.925 6.265 316.055 ;
		RECT	6.605 315.925 6.655 316.055 ;
		RECT	7.265 315.925 7.315 316.055 ;
		RECT	8.96 315.925 9.01 316.055 ;
		RECT	9.31 315.925 9.36 316.055 ;
		RECT	12.095 315.925 12.145 316.055 ;
		RECT	12.355 315.925 12.405 316.055 ;
		RECT	13.06 315.925 13.11 316.055 ;
		RECT	14.52 315.925 14.57 316.055 ;
		RECT	14.87 238.395 14.92 238.525 ;
		RECT	6.76 238.855 6.81 238.985 ;
		RECT	8.04 238.855 8.09 238.985 ;
		RECT	9.58 238.855 9.63 238.985 ;
		RECT	9.855 238.855 9.905 238.985 ;
		RECT	10.26 238.855 10.31 238.985 ;
		RECT	11.565 238.855 11.615 238.985 ;
		RECT	13.33 238.855 13.38 238.985 ;
		RECT	14.23 238.855 14.28 238.985 ;
		RECT	14.23 240.585 14.28 240.715 ;
		RECT	14.87 240.815 14.92 240.945 ;
		RECT	6.215 241.045 6.265 241.175 ;
		RECT	6.605 241.045 6.655 241.175 ;
		RECT	7.265 241.045 7.315 241.175 ;
		RECT	8.96 241.045 9.01 241.175 ;
		RECT	9.31 241.045 9.36 241.175 ;
		RECT	12.095 241.045 12.145 241.175 ;
		RECT	12.355 241.045 12.405 241.175 ;
		RECT	13.06 241.045 13.11 241.175 ;
		RECT	14.52 241.045 14.57 241.175 ;
		RECT	14.87 316.155 14.92 316.285 ;
		RECT	6.76 316.615 6.81 316.745 ;
		RECT	8.04 316.615 8.09 316.745 ;
		RECT	9.58 316.615 9.63 316.745 ;
		RECT	9.855 316.615 9.905 316.745 ;
		RECT	10.26 316.615 10.31 316.745 ;
		RECT	11.565 316.615 11.615 316.745 ;
		RECT	13.33 316.615 13.38 316.745 ;
		RECT	14.23 316.615 14.28 316.745 ;
		RECT	14.23 318.345 14.28 318.475 ;
		RECT	14.87 318.575 14.92 318.705 ;
		RECT	6.215 318.805 6.265 318.935 ;
		RECT	6.605 318.805 6.655 318.935 ;
		RECT	7.265 318.805 7.315 318.935 ;
		RECT	8.96 318.805 9.01 318.935 ;
		RECT	9.31 318.805 9.36 318.935 ;
		RECT	12.095 318.805 12.145 318.935 ;
		RECT	12.355 318.805 12.405 318.935 ;
		RECT	13.06 318.805 13.11 318.935 ;
		RECT	14.52 318.805 14.57 318.935 ;
		RECT	14.87 319.035 14.92 319.165 ;
		RECT	6.76 319.495 6.81 319.625 ;
		RECT	8.04 319.495 8.09 319.625 ;
		RECT	9.58 319.495 9.63 319.625 ;
		RECT	9.855 319.495 9.905 319.625 ;
		RECT	10.26 319.495 10.31 319.625 ;
		RECT	11.565 319.495 11.615 319.625 ;
		RECT	13.33 319.495 13.38 319.625 ;
		RECT	14.23 319.495 14.28 319.625 ;
		RECT	14.23 321.225 14.28 321.355 ;
		RECT	14.87 321.455 14.92 321.585 ;
		RECT	6.215 321.685 6.265 321.815 ;
		RECT	6.605 321.685 6.655 321.815 ;
		RECT	7.265 321.685 7.315 321.815 ;
		RECT	8.96 321.685 9.01 321.815 ;
		RECT	9.31 321.685 9.36 321.815 ;
		RECT	12.095 321.685 12.145 321.815 ;
		RECT	12.355 321.685 12.405 321.815 ;
		RECT	13.06 321.685 13.11 321.815 ;
		RECT	14.52 321.685 14.57 321.815 ;
		RECT	14.87 321.915 14.92 322.045 ;
		RECT	6.76 322.375 6.81 322.505 ;
		RECT	8.04 322.375 8.09 322.505 ;
		RECT	9.58 322.375 9.63 322.505 ;
		RECT	9.855 322.375 9.905 322.505 ;
		RECT	10.26 322.375 10.31 322.505 ;
		RECT	11.565 322.375 11.615 322.505 ;
		RECT	13.33 322.375 13.38 322.505 ;
		RECT	14.23 322.375 14.28 322.505 ;
		RECT	14.23 324.105 14.28 324.235 ;
		RECT	14.87 324.335 14.92 324.465 ;
		RECT	6.215 324.565 6.265 324.695 ;
		RECT	6.605 324.565 6.655 324.695 ;
		RECT	7.265 324.565 7.315 324.695 ;
		RECT	8.96 324.565 9.01 324.695 ;
		RECT	9.31 324.565 9.36 324.695 ;
		RECT	12.095 324.565 12.145 324.695 ;
		RECT	12.355 324.565 12.405 324.695 ;
		RECT	13.06 324.565 13.11 324.695 ;
		RECT	14.52 324.565 14.57 324.695 ;
		RECT	14.87 324.795 14.92 324.925 ;
		RECT	6.76 325.255 6.81 325.385 ;
		RECT	8.04 325.255 8.09 325.385 ;
		RECT	9.58 325.255 9.63 325.385 ;
		RECT	9.855 325.255 9.905 325.385 ;
		RECT	10.26 325.255 10.31 325.385 ;
		RECT	11.565 325.255 11.615 325.385 ;
		RECT	13.33 325.255 13.38 325.385 ;
		RECT	14.23 325.255 14.28 325.385 ;
		RECT	14.23 326.985 14.28 327.115 ;
		RECT	14.87 327.215 14.92 327.345 ;
		RECT	6.215 327.445 6.265 327.575 ;
		RECT	6.605 327.445 6.655 327.575 ;
		RECT	7.265 327.445 7.315 327.575 ;
		RECT	8.96 327.445 9.01 327.575 ;
		RECT	9.31 327.445 9.36 327.575 ;
		RECT	12.095 327.445 12.145 327.575 ;
		RECT	12.355 327.445 12.405 327.575 ;
		RECT	13.06 327.445 13.11 327.575 ;
		RECT	14.52 327.445 14.57 327.575 ;
		RECT	14.87 327.675 14.92 327.805 ;
		RECT	6.76 328.135 6.81 328.265 ;
		RECT	8.04 328.135 8.09 328.265 ;
		RECT	9.58 328.135 9.63 328.265 ;
		RECT	9.855 328.135 9.905 328.265 ;
		RECT	10.26 328.135 10.31 328.265 ;
		RECT	11.565 328.135 11.615 328.265 ;
		RECT	13.33 328.135 13.38 328.265 ;
		RECT	14.23 328.135 14.28 328.265 ;
		RECT	14.23 329.865 14.28 329.995 ;
		RECT	14.87 330.095 14.92 330.225 ;
		RECT	6.215 330.325 6.265 330.455 ;
		RECT	6.605 330.325 6.655 330.455 ;
		RECT	7.265 330.325 7.315 330.455 ;
		RECT	8.96 330.325 9.01 330.455 ;
		RECT	9.31 330.325 9.36 330.455 ;
		RECT	12.095 330.325 12.145 330.455 ;
		RECT	12.355 330.325 12.405 330.455 ;
		RECT	13.06 330.325 13.11 330.455 ;
		RECT	14.52 330.325 14.57 330.455 ;
		RECT	14.87 330.555 14.92 330.685 ;
		RECT	6.76 331.015 6.81 331.145 ;
		RECT	8.04 331.015 8.09 331.145 ;
		RECT	9.58 331.015 9.63 331.145 ;
		RECT	9.855 331.015 9.905 331.145 ;
		RECT	10.26 331.015 10.31 331.145 ;
		RECT	11.565 331.015 11.615 331.145 ;
		RECT	13.33 331.015 13.38 331.145 ;
		RECT	14.23 331.015 14.28 331.145 ;
		RECT	14.23 332.745 14.28 332.875 ;
		RECT	14.87 332.975 14.92 333.105 ;
		RECT	6.215 333.205 6.265 333.335 ;
		RECT	6.605 333.205 6.655 333.335 ;
		RECT	7.265 333.205 7.315 333.335 ;
		RECT	8.96 333.205 9.01 333.335 ;
		RECT	9.31 333.205 9.36 333.335 ;
		RECT	12.095 333.205 12.145 333.335 ;
		RECT	12.355 333.205 12.405 333.335 ;
		RECT	13.06 333.205 13.11 333.335 ;
		RECT	14.52 333.205 14.57 333.335 ;
		RECT	14.87 333.435 14.92 333.565 ;
		RECT	6.76 333.895 6.81 334.025 ;
		RECT	8.04 333.895 8.09 334.025 ;
		RECT	9.58 333.895 9.63 334.025 ;
		RECT	9.855 333.895 9.905 334.025 ;
		RECT	10.26 333.895 10.31 334.025 ;
		RECT	11.565 333.895 11.615 334.025 ;
		RECT	13.33 333.895 13.38 334.025 ;
		RECT	14.23 333.895 14.28 334.025 ;
		RECT	14.23 335.625 14.28 335.755 ;
		RECT	14.87 335.855 14.92 335.985 ;
		RECT	6.215 336.085 6.265 336.215 ;
		RECT	6.605 336.085 6.655 336.215 ;
		RECT	7.265 336.085 7.315 336.215 ;
		RECT	8.96 336.085 9.01 336.215 ;
		RECT	9.31 336.085 9.36 336.215 ;
		RECT	12.095 336.085 12.145 336.215 ;
		RECT	12.355 336.085 12.405 336.215 ;
		RECT	13.06 336.085 13.11 336.215 ;
		RECT	14.52 336.085 14.57 336.215 ;
		RECT	14.87 336.315 14.92 336.445 ;
		RECT	6.76 336.775 6.81 336.905 ;
		RECT	8.04 336.775 8.09 336.905 ;
		RECT	9.58 336.775 9.63 336.905 ;
		RECT	9.855 336.775 9.905 336.905 ;
		RECT	10.26 336.775 10.31 336.905 ;
		RECT	11.565 336.775 11.615 336.905 ;
		RECT	13.33 336.775 13.38 336.905 ;
		RECT	14.23 336.775 14.28 336.905 ;
		RECT	14.23 338.505 14.28 338.635 ;
		RECT	14.87 338.735 14.92 338.865 ;
		RECT	6.215 338.965 6.265 339.095 ;
		RECT	6.605 338.965 6.655 339.095 ;
		RECT	7.265 338.965 7.315 339.095 ;
		RECT	8.96 338.965 9.01 339.095 ;
		RECT	9.31 338.965 9.36 339.095 ;
		RECT	12.095 338.965 12.145 339.095 ;
		RECT	12.355 338.965 12.405 339.095 ;
		RECT	13.06 338.965 13.11 339.095 ;
		RECT	14.52 338.965 14.57 339.095 ;
		RECT	14.87 339.195 14.92 339.325 ;
		RECT	6.76 339.655 6.81 339.785 ;
		RECT	8.04 339.655 8.09 339.785 ;
		RECT	9.58 339.655 9.63 339.785 ;
		RECT	9.855 339.655 9.905 339.785 ;
		RECT	10.26 339.655 10.31 339.785 ;
		RECT	11.565 339.655 11.615 339.785 ;
		RECT	13.33 339.655 13.38 339.785 ;
		RECT	14.23 339.655 14.28 339.785 ;
		RECT	14.23 341.385 14.28 341.515 ;
		RECT	14.87 341.615 14.92 341.745 ;
		RECT	6.215 341.845 6.265 341.975 ;
		RECT	6.605 341.845 6.655 341.975 ;
		RECT	7.265 341.845 7.315 341.975 ;
		RECT	8.96 341.845 9.01 341.975 ;
		RECT	9.31 341.845 9.36 341.975 ;
		RECT	12.095 341.845 12.145 341.975 ;
		RECT	12.355 341.845 12.405 341.975 ;
		RECT	13.06 341.845 13.11 341.975 ;
		RECT	14.52 341.845 14.57 341.975 ;
		RECT	14.87 342.075 14.92 342.205 ;
		RECT	6.76 342.535 6.81 342.665 ;
		RECT	8.04 342.535 8.09 342.665 ;
		RECT	9.58 342.535 9.63 342.665 ;
		RECT	9.855 342.535 9.905 342.665 ;
		RECT	10.26 342.535 10.31 342.665 ;
		RECT	11.565 342.535 11.615 342.665 ;
		RECT	13.33 342.535 13.38 342.665 ;
		RECT	14.23 342.535 14.28 342.665 ;
		RECT	14.23 344.265 14.28 344.395 ;
		RECT	14.87 344.495 14.92 344.625 ;
		RECT	6.215 344.725 6.265 344.855 ;
		RECT	6.605 344.725 6.655 344.855 ;
		RECT	7.265 344.725 7.315 344.855 ;
		RECT	8.96 344.725 9.01 344.855 ;
		RECT	9.31 344.725 9.36 344.855 ;
		RECT	12.095 344.725 12.145 344.855 ;
		RECT	12.355 344.725 12.405 344.855 ;
		RECT	13.06 344.725 13.11 344.855 ;
		RECT	14.52 344.725 14.57 344.855 ;
		RECT	14.87 241.275 14.92 241.405 ;
		RECT	6.76 241.735 6.81 241.865 ;
		RECT	8.04 241.735 8.09 241.865 ;
		RECT	9.58 241.735 9.63 241.865 ;
		RECT	9.855 241.735 9.905 241.865 ;
		RECT	10.26 241.735 10.31 241.865 ;
		RECT	11.565 241.735 11.615 241.865 ;
		RECT	13.33 241.735 13.38 241.865 ;
		RECT	14.23 241.735 14.28 241.865 ;
		RECT	14.23 243.465 14.28 243.595 ;
		RECT	14.87 243.695 14.92 243.825 ;
		RECT	6.215 243.925 6.265 244.055 ;
		RECT	6.605 243.925 6.655 244.055 ;
		RECT	7.265 243.925 7.315 244.055 ;
		RECT	8.96 243.925 9.01 244.055 ;
		RECT	9.31 243.925 9.36 244.055 ;
		RECT	12.095 243.925 12.145 244.055 ;
		RECT	12.355 243.925 12.405 244.055 ;
		RECT	13.06 243.925 13.11 244.055 ;
		RECT	14.52 243.925 14.57 244.055 ;
		RECT	14.87 344.955 14.92 345.085 ;
		RECT	6.76 345.415 6.81 345.545 ;
		RECT	8.04 345.415 8.09 345.545 ;
		RECT	9.58 345.415 9.63 345.545 ;
		RECT	9.855 345.415 9.905 345.545 ;
		RECT	10.26 345.415 10.31 345.545 ;
		RECT	11.565 345.415 11.615 345.545 ;
		RECT	13.33 345.415 13.38 345.545 ;
		RECT	14.23 345.415 14.28 345.545 ;
		RECT	14.23 347.145 14.28 347.275 ;
		RECT	14.87 347.375 14.92 347.505 ;
		RECT	6.215 347.605 6.265 347.735 ;
		RECT	6.605 347.605 6.655 347.735 ;
		RECT	7.265 347.605 7.315 347.735 ;
		RECT	8.96 347.605 9.01 347.735 ;
		RECT	9.31 347.605 9.36 347.735 ;
		RECT	12.095 347.605 12.145 347.735 ;
		RECT	12.355 347.605 12.405 347.735 ;
		RECT	13.06 347.605 13.11 347.735 ;
		RECT	14.52 347.605 14.57 347.735 ;
		RECT	14.87 347.835 14.92 347.965 ;
		RECT	6.76 348.295 6.81 348.425 ;
		RECT	8.04 348.295 8.09 348.425 ;
		RECT	9.58 348.295 9.63 348.425 ;
		RECT	9.855 348.295 9.905 348.425 ;
		RECT	10.26 348.295 10.31 348.425 ;
		RECT	11.565 348.295 11.615 348.425 ;
		RECT	13.33 348.295 13.38 348.425 ;
		RECT	14.23 348.295 14.28 348.425 ;
		RECT	14.23 350.025 14.28 350.155 ;
		RECT	14.87 350.255 14.92 350.385 ;
		RECT	6.215 350.485 6.265 350.615 ;
		RECT	6.605 350.485 6.655 350.615 ;
		RECT	7.265 350.485 7.315 350.615 ;
		RECT	8.96 350.485 9.01 350.615 ;
		RECT	9.31 350.485 9.36 350.615 ;
		RECT	12.095 350.485 12.145 350.615 ;
		RECT	12.355 350.485 12.405 350.615 ;
		RECT	13.06 350.485 13.11 350.615 ;
		RECT	14.52 350.485 14.57 350.615 ;
		RECT	14.87 350.715 14.92 350.845 ;
		RECT	6.76 351.175 6.81 351.305 ;
		RECT	8.04 351.175 8.09 351.305 ;
		RECT	9.58 351.175 9.63 351.305 ;
		RECT	9.855 351.175 9.905 351.305 ;
		RECT	10.26 351.175 10.31 351.305 ;
		RECT	11.565 351.175 11.615 351.305 ;
		RECT	13.33 351.175 13.38 351.305 ;
		RECT	14.23 351.175 14.28 351.305 ;
		RECT	14.23 352.905 14.28 353.035 ;
		RECT	14.87 353.135 14.92 353.265 ;
		RECT	6.215 353.365 6.265 353.495 ;
		RECT	6.605 353.365 6.655 353.495 ;
		RECT	7.265 353.365 7.315 353.495 ;
		RECT	8.96 353.365 9.01 353.495 ;
		RECT	9.31 353.365 9.36 353.495 ;
		RECT	12.095 353.365 12.145 353.495 ;
		RECT	12.355 353.365 12.405 353.495 ;
		RECT	13.06 353.365 13.11 353.495 ;
		RECT	14.52 353.365 14.57 353.495 ;
		RECT	14.87 353.595 14.92 353.725 ;
		RECT	6.76 354.055 6.81 354.185 ;
		RECT	8.04 354.055 8.09 354.185 ;
		RECT	9.58 354.055 9.63 354.185 ;
		RECT	9.855 354.055 9.905 354.185 ;
		RECT	10.26 354.055 10.31 354.185 ;
		RECT	11.565 354.055 11.615 354.185 ;
		RECT	13.33 354.055 13.38 354.185 ;
		RECT	14.23 354.055 14.28 354.185 ;
		RECT	14.23 355.785 14.28 355.915 ;
		RECT	14.87 356.015 14.92 356.145 ;
		RECT	6.215 356.245 6.265 356.375 ;
		RECT	6.605 356.245 6.655 356.375 ;
		RECT	7.265 356.245 7.315 356.375 ;
		RECT	8.96 356.245 9.01 356.375 ;
		RECT	9.31 356.245 9.36 356.375 ;
		RECT	12.095 356.245 12.145 356.375 ;
		RECT	12.355 356.245 12.405 356.375 ;
		RECT	13.06 356.245 13.11 356.375 ;
		RECT	14.52 356.245 14.57 356.375 ;
		RECT	14.87 356.475 14.92 356.605 ;
		RECT	6.76 356.935 6.81 357.065 ;
		RECT	8.04 356.935 8.09 357.065 ;
		RECT	9.58 356.935 9.63 357.065 ;
		RECT	9.855 356.935 9.905 357.065 ;
		RECT	10.26 356.935 10.31 357.065 ;
		RECT	11.565 356.935 11.615 357.065 ;
		RECT	13.33 356.935 13.38 357.065 ;
		RECT	14.23 356.935 14.28 357.065 ;
		RECT	14.23 358.665 14.28 358.795 ;
		RECT	14.87 358.895 14.92 359.025 ;
		RECT	6.215 359.125 6.265 359.255 ;
		RECT	6.605 359.125 6.655 359.255 ;
		RECT	7.265 359.125 7.315 359.255 ;
		RECT	8.96 359.125 9.01 359.255 ;
		RECT	9.31 359.125 9.36 359.255 ;
		RECT	12.095 359.125 12.145 359.255 ;
		RECT	12.355 359.125 12.405 359.255 ;
		RECT	13.06 359.125 13.11 359.255 ;
		RECT	14.52 359.125 14.57 359.255 ;
		RECT	14.87 359.355 14.92 359.485 ;
		RECT	6.76 359.815 6.81 359.945 ;
		RECT	8.04 359.815 8.09 359.945 ;
		RECT	9.58 359.815 9.63 359.945 ;
		RECT	9.855 359.815 9.905 359.945 ;
		RECT	10.26 359.815 10.31 359.945 ;
		RECT	11.565 359.815 11.615 359.945 ;
		RECT	13.33 359.815 13.38 359.945 ;
		RECT	14.23 359.815 14.28 359.945 ;
		RECT	14.23 361.545 14.28 361.675 ;
		RECT	14.87 361.775 14.92 361.905 ;
		RECT	6.215 362.005 6.265 362.135 ;
		RECT	6.605 362.005 6.655 362.135 ;
		RECT	7.265 362.005 7.315 362.135 ;
		RECT	8.96 362.005 9.01 362.135 ;
		RECT	9.31 362.005 9.36 362.135 ;
		RECT	12.095 362.005 12.145 362.135 ;
		RECT	12.355 362.005 12.405 362.135 ;
		RECT	13.06 362.005 13.11 362.135 ;
		RECT	14.52 362.005 14.57 362.135 ;
		RECT	14.87 362.235 14.92 362.365 ;
		RECT	6.76 362.695 6.81 362.825 ;
		RECT	8.04 362.695 8.09 362.825 ;
		RECT	9.58 362.695 9.63 362.825 ;
		RECT	9.855 362.695 9.905 362.825 ;
		RECT	10.26 362.695 10.31 362.825 ;
		RECT	11.565 362.695 11.615 362.825 ;
		RECT	13.33 362.695 13.38 362.825 ;
		RECT	14.23 362.695 14.28 362.825 ;
		RECT	14.23 364.425 14.28 364.555 ;
		RECT	14.87 364.655 14.92 364.785 ;
		RECT	6.215 364.885 6.265 365.015 ;
		RECT	6.605 364.885 6.655 365.015 ;
		RECT	7.265 364.885 7.315 365.015 ;
		RECT	8.96 364.885 9.01 365.015 ;
		RECT	9.31 364.885 9.36 365.015 ;
		RECT	12.095 364.885 12.145 365.015 ;
		RECT	12.355 364.885 12.405 365.015 ;
		RECT	13.06 364.885 13.11 365.015 ;
		RECT	14.52 364.885 14.57 365.015 ;
		RECT	14.87 365.115 14.92 365.245 ;
		RECT	6.76 365.575 6.81 365.705 ;
		RECT	8.04 365.575 8.09 365.705 ;
		RECT	9.58 365.575 9.63 365.705 ;
		RECT	9.855 365.575 9.905 365.705 ;
		RECT	10.26 365.575 10.31 365.705 ;
		RECT	11.565 365.575 11.615 365.705 ;
		RECT	13.33 365.575 13.38 365.705 ;
		RECT	14.23 365.575 14.28 365.705 ;
		RECT	14.23 367.305 14.28 367.435 ;
		RECT	14.87 367.535 14.92 367.665 ;
		RECT	6.215 367.765 6.265 367.895 ;
		RECT	6.605 367.765 6.655 367.895 ;
		RECT	7.265 367.765 7.315 367.895 ;
		RECT	8.96 367.765 9.01 367.895 ;
		RECT	9.31 367.765 9.36 367.895 ;
		RECT	12.095 367.765 12.145 367.895 ;
		RECT	12.355 367.765 12.405 367.895 ;
		RECT	13.06 367.765 13.11 367.895 ;
		RECT	14.52 367.765 14.57 367.895 ;
		RECT	14.87 367.995 14.92 368.125 ;
		RECT	6.76 368.455 6.81 368.585 ;
		RECT	8.04 368.455 8.09 368.585 ;
		RECT	9.58 368.455 9.63 368.585 ;
		RECT	9.855 368.455 9.905 368.585 ;
		RECT	10.26 368.455 10.31 368.585 ;
		RECT	11.565 368.455 11.615 368.585 ;
		RECT	13.33 368.455 13.38 368.585 ;
		RECT	14.23 368.455 14.28 368.585 ;
		RECT	14.23 370.185 14.28 370.315 ;
		RECT	14.87 370.415 14.92 370.545 ;
		RECT	6.215 370.645 6.265 370.775 ;
		RECT	6.605 370.645 6.655 370.775 ;
		RECT	7.265 370.645 7.315 370.775 ;
		RECT	8.96 370.645 9.01 370.775 ;
		RECT	9.31 370.645 9.36 370.775 ;
		RECT	12.095 370.645 12.145 370.775 ;
		RECT	12.355 370.645 12.405 370.775 ;
		RECT	13.06 370.645 13.11 370.775 ;
		RECT	14.52 370.645 14.57 370.775 ;
		RECT	14.87 370.875 14.92 371.005 ;
		RECT	6.76 371.335 6.81 371.465 ;
		RECT	8.04 371.335 8.09 371.465 ;
		RECT	9.58 371.335 9.63 371.465 ;
		RECT	9.855 371.335 9.905 371.465 ;
		RECT	10.26 371.335 10.31 371.465 ;
		RECT	11.565 371.335 11.615 371.465 ;
		RECT	13.33 371.335 13.38 371.465 ;
		RECT	14.23 371.335 14.28 371.465 ;
		RECT	14.23 373.065 14.28 373.195 ;
		RECT	14.87 373.295 14.92 373.425 ;
		RECT	6.215 373.525 6.265 373.655 ;
		RECT	6.605 373.525 6.655 373.655 ;
		RECT	7.265 373.525 7.315 373.655 ;
		RECT	8.96 373.525 9.01 373.655 ;
		RECT	9.31 373.525 9.36 373.655 ;
		RECT	12.095 373.525 12.145 373.655 ;
		RECT	12.355 373.525 12.405 373.655 ;
		RECT	13.06 373.525 13.11 373.655 ;
		RECT	14.52 373.525 14.57 373.655 ;
		RECT	14.87 244.155 14.92 244.285 ;
		RECT	6.76 244.615 6.81 244.745 ;
		RECT	8.04 244.615 8.09 244.745 ;
		RECT	9.58 244.615 9.63 244.745 ;
		RECT	9.855 244.615 9.905 244.745 ;
		RECT	10.26 244.615 10.31 244.745 ;
		RECT	11.565 244.615 11.615 244.745 ;
		RECT	13.33 244.615 13.38 244.745 ;
		RECT	14.23 244.615 14.28 244.745 ;
		RECT	14.23 246.345 14.28 246.475 ;
		RECT	14.87 246.575 14.92 246.705 ;
		RECT	6.215 246.805 6.265 246.935 ;
		RECT	6.605 246.805 6.655 246.935 ;
		RECT	7.265 246.805 7.315 246.935 ;
		RECT	8.96 246.805 9.01 246.935 ;
		RECT	9.31 246.805 9.36 246.935 ;
		RECT	12.095 246.805 12.145 246.935 ;
		RECT	12.355 246.805 12.405 246.935 ;
		RECT	13.06 246.805 13.11 246.935 ;
		RECT	14.52 246.805 14.57 246.935 ;
		RECT	14.87 373.755 14.92 373.885 ;
		RECT	6.76 374.215 6.81 374.345 ;
		RECT	8.04 374.215 8.09 374.345 ;
		RECT	9.58 374.215 9.63 374.345 ;
		RECT	9.855 374.215 9.905 374.345 ;
		RECT	10.26 374.215 10.31 374.345 ;
		RECT	11.565 374.215 11.615 374.345 ;
		RECT	13.33 374.215 13.38 374.345 ;
		RECT	14.23 374.215 14.28 374.345 ;
		RECT	14.23 375.945 14.28 376.075 ;
		RECT	14.87 376.175 14.92 376.305 ;
		RECT	6.215 376.405 6.265 376.535 ;
		RECT	6.605 376.405 6.655 376.535 ;
		RECT	7.265 376.405 7.315 376.535 ;
		RECT	8.96 376.405 9.01 376.535 ;
		RECT	9.31 376.405 9.36 376.535 ;
		RECT	12.095 376.405 12.145 376.535 ;
		RECT	12.355 376.405 12.405 376.535 ;
		RECT	13.06 376.405 13.11 376.535 ;
		RECT	14.52 376.405 14.57 376.535 ;
		RECT	14.87 376.635 14.92 376.765 ;
		RECT	6.76 377.095 6.81 377.225 ;
		RECT	8.04 377.095 8.09 377.225 ;
		RECT	9.58 377.095 9.63 377.225 ;
		RECT	9.855 377.095 9.905 377.225 ;
		RECT	10.26 377.095 10.31 377.225 ;
		RECT	11.565 377.095 11.615 377.225 ;
		RECT	13.33 377.095 13.38 377.225 ;
		RECT	14.23 377.095 14.28 377.225 ;
		RECT	14.23 378.825 14.28 378.955 ;
		RECT	14.87 379.055 14.92 379.185 ;
		RECT	6.215 379.285 6.265 379.415 ;
		RECT	6.605 379.285 6.655 379.415 ;
		RECT	7.265 379.285 7.315 379.415 ;
		RECT	8.96 379.285 9.01 379.415 ;
		RECT	9.31 379.285 9.36 379.415 ;
		RECT	12.095 379.285 12.145 379.415 ;
		RECT	12.355 379.285 12.405 379.415 ;
		RECT	13.06 379.285 13.11 379.415 ;
		RECT	14.52 379.285 14.57 379.415 ;
		RECT	14.87 379.515 14.92 379.645 ;
		RECT	6.76 379.975 6.81 380.105 ;
		RECT	8.04 379.975 8.09 380.105 ;
		RECT	9.58 379.975 9.63 380.105 ;
		RECT	9.855 379.975 9.905 380.105 ;
		RECT	10.26 379.975 10.31 380.105 ;
		RECT	11.565 379.975 11.615 380.105 ;
		RECT	13.33 379.975 13.38 380.105 ;
		RECT	14.23 379.975 14.28 380.105 ;
		RECT	14.23 381.705 14.28 381.835 ;
		RECT	14.87 381.935 14.92 382.065 ;
		RECT	6.215 382.165 6.265 382.295 ;
		RECT	6.605 382.165 6.655 382.295 ;
		RECT	7.265 382.165 7.315 382.295 ;
		RECT	8.96 382.165 9.01 382.295 ;
		RECT	9.31 382.165 9.36 382.295 ;
		RECT	12.095 382.165 12.145 382.295 ;
		RECT	12.355 382.165 12.405 382.295 ;
		RECT	13.06 382.165 13.11 382.295 ;
		RECT	14.52 382.165 14.57 382.295 ;
		RECT	14.87 382.395 14.92 382.525 ;
		RECT	6.76 382.855 6.81 382.985 ;
		RECT	8.04 382.855 8.09 382.985 ;
		RECT	9.58 382.855 9.63 382.985 ;
		RECT	9.855 382.855 9.905 382.985 ;
		RECT	10.26 382.855 10.31 382.985 ;
		RECT	11.565 382.855 11.615 382.985 ;
		RECT	13.33 382.855 13.38 382.985 ;
		RECT	14.23 382.855 14.28 382.985 ;
		RECT	14.23 384.585 14.28 384.715 ;
		RECT	14.87 384.815 14.92 384.945 ;
		RECT	6.215 385.045 6.265 385.175 ;
		RECT	6.605 385.045 6.655 385.175 ;
		RECT	7.265 385.045 7.315 385.175 ;
		RECT	8.96 385.045 9.01 385.175 ;
		RECT	9.31 385.045 9.36 385.175 ;
		RECT	12.095 385.045 12.145 385.175 ;
		RECT	12.355 385.045 12.405 385.175 ;
		RECT	13.06 385.045 13.11 385.175 ;
		RECT	14.52 385.045 14.57 385.175 ;
		RECT	14.87 385.275 14.92 385.405 ;
		RECT	6.76 385.735 6.81 385.865 ;
		RECT	8.04 385.735 8.09 385.865 ;
		RECT	9.58 385.735 9.63 385.865 ;
		RECT	9.855 385.735 9.905 385.865 ;
		RECT	10.26 385.735 10.31 385.865 ;
		RECT	11.565 385.735 11.615 385.865 ;
		RECT	13.33 385.735 13.38 385.865 ;
		RECT	14.23 385.735 14.28 385.865 ;
		RECT	14.23 387.465 14.28 387.595 ;
		RECT	14.87 387.695 14.92 387.825 ;
		RECT	6.215 387.925 6.265 388.055 ;
		RECT	6.605 387.925 6.655 388.055 ;
		RECT	7.265 387.925 7.315 388.055 ;
		RECT	8.96 387.925 9.01 388.055 ;
		RECT	9.31 387.925 9.36 388.055 ;
		RECT	12.095 387.925 12.145 388.055 ;
		RECT	12.355 387.925 12.405 388.055 ;
		RECT	13.06 387.925 13.11 388.055 ;
		RECT	14.52 387.925 14.57 388.055 ;
		RECT	14.87 388.155 14.92 388.285 ;
		RECT	6.76 388.615 6.81 388.745 ;
		RECT	8.04 388.615 8.09 388.745 ;
		RECT	9.58 388.615 9.63 388.745 ;
		RECT	9.855 388.615 9.905 388.745 ;
		RECT	10.26 388.615 10.31 388.745 ;
		RECT	11.565 388.615 11.615 388.745 ;
		RECT	13.33 388.615 13.38 388.745 ;
		RECT	14.23 388.615 14.28 388.745 ;
		RECT	14.23 390.345 14.28 390.475 ;
		RECT	14.87 390.575 14.92 390.705 ;
		RECT	6.215 390.805 6.265 390.935 ;
		RECT	6.605 390.805 6.655 390.935 ;
		RECT	7.265 390.805 7.315 390.935 ;
		RECT	8.96 390.805 9.01 390.935 ;
		RECT	9.31 390.805 9.36 390.935 ;
		RECT	12.095 390.805 12.145 390.935 ;
		RECT	12.355 390.805 12.405 390.935 ;
		RECT	13.06 390.805 13.11 390.935 ;
		RECT	14.52 390.805 14.57 390.935 ;
		RECT	14.87 391.035 14.92 391.165 ;
		RECT	6.76 391.495 6.81 391.625 ;
		RECT	8.04 391.495 8.09 391.625 ;
		RECT	9.58 391.495 9.63 391.625 ;
		RECT	9.855 391.495 9.905 391.625 ;
		RECT	10.26 391.495 10.31 391.625 ;
		RECT	11.565 391.495 11.615 391.625 ;
		RECT	13.33 391.495 13.38 391.625 ;
		RECT	14.23 391.495 14.28 391.625 ;
		RECT	14.23 393.225 14.28 393.355 ;
		RECT	14.87 393.455 14.92 393.585 ;
		RECT	6.215 393.685 6.265 393.815 ;
		RECT	6.605 393.685 6.655 393.815 ;
		RECT	7.265 393.685 7.315 393.815 ;
		RECT	8.96 393.685 9.01 393.815 ;
		RECT	9.31 393.685 9.36 393.815 ;
		RECT	12.095 393.685 12.145 393.815 ;
		RECT	12.355 393.685 12.405 393.815 ;
		RECT	13.06 393.685 13.11 393.815 ;
		RECT	14.52 393.685 14.57 393.815 ;
		RECT	14.87 393.915 14.92 394.045 ;
		RECT	6.76 394.375 6.81 394.505 ;
		RECT	8.04 394.375 8.09 394.505 ;
		RECT	9.58 394.375 9.63 394.505 ;
		RECT	9.855 394.375 9.905 394.505 ;
		RECT	10.26 394.375 10.31 394.505 ;
		RECT	11.565 394.375 11.615 394.505 ;
		RECT	13.33 394.375 13.38 394.505 ;
		RECT	14.23 394.375 14.28 394.505 ;
		RECT	14.23 396.105 14.28 396.235 ;
		RECT	14.87 396.335 14.92 396.465 ;
		RECT	6.215 396.565 6.265 396.695 ;
		RECT	6.605 396.565 6.655 396.695 ;
		RECT	7.265 396.565 7.315 396.695 ;
		RECT	8.96 396.565 9.01 396.695 ;
		RECT	9.31 396.565 9.36 396.695 ;
		RECT	12.095 396.565 12.145 396.695 ;
		RECT	12.355 396.565 12.405 396.695 ;
		RECT	13.06 396.565 13.11 396.695 ;
		RECT	14.52 396.565 14.57 396.695 ;
		RECT	14.87 396.795 14.92 396.925 ;
		RECT	6.76 397.255 6.81 397.385 ;
		RECT	8.04 397.255 8.09 397.385 ;
		RECT	9.58 397.255 9.63 397.385 ;
		RECT	9.855 397.255 9.905 397.385 ;
		RECT	10.26 397.255 10.31 397.385 ;
		RECT	11.565 397.255 11.615 397.385 ;
		RECT	13.33 397.255 13.38 397.385 ;
		RECT	14.23 397.255 14.28 397.385 ;
		RECT	14.23 398.985 14.28 399.115 ;
		RECT	14.87 399.215 14.92 399.345 ;
		RECT	6.215 399.445 6.265 399.575 ;
		RECT	6.605 399.445 6.655 399.575 ;
		RECT	7.265 399.445 7.315 399.575 ;
		RECT	8.96 399.445 9.01 399.575 ;
		RECT	9.31 399.445 9.36 399.575 ;
		RECT	12.095 399.445 12.145 399.575 ;
		RECT	12.355 399.445 12.405 399.575 ;
		RECT	13.06 399.445 13.11 399.575 ;
		RECT	14.52 399.445 14.57 399.575 ;
		RECT	14.87 399.675 14.92 399.805 ;
		RECT	6.76 400.135 6.81 400.265 ;
		RECT	8.04 400.135 8.09 400.265 ;
		RECT	9.58 400.135 9.63 400.265 ;
		RECT	9.855 400.135 9.905 400.265 ;
		RECT	10.26 400.135 10.31 400.265 ;
		RECT	11.565 400.135 11.615 400.265 ;
		RECT	13.33 400.135 13.38 400.265 ;
		RECT	14.23 400.135 14.28 400.265 ;
		RECT	14.23 401.865 14.28 401.995 ;
		RECT	14.87 402.095 14.92 402.225 ;
		RECT	6.215 402.325 6.265 402.455 ;
		RECT	6.605 402.325 6.655 402.455 ;
		RECT	7.265 402.325 7.315 402.455 ;
		RECT	8.96 402.325 9.01 402.455 ;
		RECT	9.31 402.325 9.36 402.455 ;
		RECT	12.095 402.325 12.145 402.455 ;
		RECT	12.355 402.325 12.405 402.455 ;
		RECT	13.06 402.325 13.11 402.455 ;
		RECT	14.52 402.325 14.57 402.455 ;
		RECT	14.87 247.035 14.92 247.165 ;
		RECT	6.76 247.495 6.81 247.625 ;
		RECT	8.04 247.495 8.09 247.625 ;
		RECT	9.58 247.495 9.63 247.625 ;
		RECT	9.855 247.495 9.905 247.625 ;
		RECT	10.26 247.495 10.31 247.625 ;
		RECT	11.565 247.495 11.615 247.625 ;
		RECT	13.33 247.495 13.38 247.625 ;
		RECT	14.23 247.495 14.28 247.625 ;
		RECT	14.23 249.225 14.28 249.355 ;
		RECT	14.87 249.455 14.92 249.585 ;
		RECT	6.215 249.685 6.265 249.815 ;
		RECT	6.605 249.685 6.655 249.815 ;
		RECT	7.265 249.685 7.315 249.815 ;
		RECT	8.96 249.685 9.01 249.815 ;
		RECT	9.31 249.685 9.36 249.815 ;
		RECT	12.095 249.685 12.145 249.815 ;
		RECT	12.355 249.685 12.405 249.815 ;
		RECT	13.06 249.685 13.11 249.815 ;
		RECT	14.52 249.685 14.57 249.815 ;
		RECT	14.87 402.555 14.92 402.685 ;
		RECT	6.76 403.015 6.81 403.145 ;
		RECT	8.04 403.015 8.09 403.145 ;
		RECT	9.58 403.015 9.63 403.145 ;
		RECT	9.855 403.015 9.905 403.145 ;
		RECT	10.26 403.015 10.31 403.145 ;
		RECT	11.565 403.015 11.615 403.145 ;
		RECT	13.33 403.015 13.38 403.145 ;
		RECT	14.23 403.015 14.28 403.145 ;
		RECT	14.23 404.745 14.28 404.875 ;
		RECT	14.87 404.975 14.92 405.105 ;
		RECT	6.215 405.205 6.265 405.335 ;
		RECT	6.605 405.205 6.655 405.335 ;
		RECT	7.265 405.205 7.315 405.335 ;
		RECT	8.96 405.205 9.01 405.335 ;
		RECT	9.31 405.205 9.36 405.335 ;
		RECT	12.095 405.205 12.145 405.335 ;
		RECT	12.355 405.205 12.405 405.335 ;
		RECT	13.06 405.205 13.11 405.335 ;
		RECT	14.52 405.205 14.57 405.335 ;
		RECT	14.87 405.435 14.92 405.565 ;
		RECT	6.76 405.895 6.81 406.025 ;
		RECT	8.04 405.895 8.09 406.025 ;
		RECT	9.58 405.895 9.63 406.025 ;
		RECT	9.855 405.895 9.905 406.025 ;
		RECT	10.26 405.895 10.31 406.025 ;
		RECT	11.565 405.895 11.615 406.025 ;
		RECT	13.33 405.895 13.38 406.025 ;
		RECT	14.23 405.895 14.28 406.025 ;
		RECT	14.23 407.625 14.28 407.755 ;
		RECT	14.87 407.855 14.92 407.985 ;
		RECT	6.215 408.085 6.265 408.215 ;
		RECT	6.605 408.085 6.655 408.215 ;
		RECT	7.265 408.085 7.315 408.215 ;
		RECT	8.96 408.085 9.01 408.215 ;
		RECT	9.31 408.085 9.36 408.215 ;
		RECT	12.095 408.085 12.145 408.215 ;
		RECT	12.355 408.085 12.405 408.215 ;
		RECT	13.06 408.085 13.11 408.215 ;
		RECT	14.52 408.085 14.57 408.215 ;
		RECT	14.87 408.315 14.92 408.445 ;
		RECT	6.76 408.775 6.81 408.905 ;
		RECT	8.04 408.775 8.09 408.905 ;
		RECT	9.58 408.775 9.63 408.905 ;
		RECT	9.855 408.775 9.905 408.905 ;
		RECT	10.26 408.775 10.31 408.905 ;
		RECT	11.565 408.775 11.615 408.905 ;
		RECT	13.33 408.775 13.38 408.905 ;
		RECT	14.23 408.775 14.28 408.905 ;
		RECT	14.23 410.505 14.28 410.635 ;
		RECT	14.87 410.735 14.92 410.865 ;
		RECT	6.215 410.965 6.265 411.095 ;
		RECT	6.605 410.965 6.655 411.095 ;
		RECT	7.265 410.965 7.315 411.095 ;
		RECT	8.96 410.965 9.01 411.095 ;
		RECT	9.31 410.965 9.36 411.095 ;
		RECT	12.095 410.965 12.145 411.095 ;
		RECT	12.355 410.965 12.405 411.095 ;
		RECT	13.06 410.965 13.11 411.095 ;
		RECT	14.52 410.965 14.57 411.095 ;
		RECT	14.87 249.915 14.92 250.045 ;
		RECT	6.76 250.375 6.81 250.505 ;
		RECT	8.04 250.375 8.09 250.505 ;
		RECT	9.58 250.375 9.63 250.505 ;
		RECT	9.855 250.375 9.905 250.505 ;
		RECT	10.26 250.375 10.31 250.505 ;
		RECT	11.565 250.375 11.615 250.505 ;
		RECT	13.33 250.375 13.38 250.505 ;
		RECT	14.23 250.375 14.28 250.505 ;
		RECT	14.23 252.105 14.28 252.235 ;
		RECT	14.87 252.335 14.92 252.465 ;
		RECT	6.215 252.565 6.265 252.695 ;
		RECT	6.605 252.565 6.655 252.695 ;
		RECT	7.265 252.565 7.315 252.695 ;
		RECT	8.96 252.565 9.01 252.695 ;
		RECT	9.31 252.565 9.36 252.695 ;
		RECT	12.095 252.565 12.145 252.695 ;
		RECT	12.355 252.565 12.405 252.695 ;
		RECT	13.06 252.565 13.11 252.695 ;
		RECT	14.52 252.565 14.57 252.695 ;
		RECT	14.87 252.795 14.92 252.925 ;
		RECT	6.76 253.255 6.81 253.385 ;
		RECT	8.04 253.255 8.09 253.385 ;
		RECT	9.58 253.255 9.63 253.385 ;
		RECT	9.855 253.255 9.905 253.385 ;
		RECT	10.26 253.255 10.31 253.385 ;
		RECT	11.565 253.255 11.615 253.385 ;
		RECT	13.33 253.255 13.38 253.385 ;
		RECT	14.23 253.255 14.28 253.385 ;
		RECT	14.23 254.985 14.28 255.115 ;
		RECT	14.87 255.215 14.92 255.345 ;
		RECT	6.215 255.445 6.265 255.575 ;
		RECT	6.605 255.445 6.655 255.575 ;
		RECT	7.265 255.445 7.315 255.575 ;
		RECT	8.96 255.445 9.01 255.575 ;
		RECT	9.31 255.445 9.36 255.575 ;
		RECT	12.095 255.445 12.145 255.575 ;
		RECT	12.355 255.445 12.405 255.575 ;
		RECT	13.06 255.445 13.11 255.575 ;
		RECT	14.52 255.445 14.57 255.575 ;
		RECT	14.87 255.675 14.92 255.805 ;
		RECT	6.76 256.135 6.81 256.265 ;
		RECT	8.04 256.135 8.09 256.265 ;
		RECT	9.58 256.135 9.63 256.265 ;
		RECT	9.855 256.135 9.905 256.265 ;
		RECT	10.26 256.135 10.31 256.265 ;
		RECT	11.565 256.135 11.615 256.265 ;
		RECT	13.33 256.135 13.38 256.265 ;
		RECT	14.23 256.135 14.28 256.265 ;
		RECT	14.23 257.865 14.28 257.995 ;
		RECT	14.87 258.095 14.92 258.225 ;
		RECT	6.215 258.325 6.265 258.455 ;
		RECT	6.605 258.325 6.655 258.455 ;
		RECT	7.265 258.325 7.315 258.455 ;
		RECT	8.96 258.325 9.01 258.455 ;
		RECT	9.31 258.325 9.36 258.455 ;
		RECT	12.095 258.325 12.145 258.455 ;
		RECT	12.355 258.325 12.405 258.455 ;
		RECT	13.06 258.325 13.11 258.455 ;
		RECT	14.52 258.325 14.57 258.455 ;
		RECT	14.87 411.195 14.92 411.325 ;
		RECT	6.76 411.655 6.81 411.785 ;
		RECT	8.04 411.655 8.09 411.785 ;
		RECT	9.58 411.655 9.63 411.785 ;
		RECT	9.855 411.655 9.905 411.785 ;
		RECT	10.26 411.655 10.31 411.785 ;
		RECT	11.565 411.655 11.615 411.785 ;
		RECT	13.33 411.655 13.38 411.785 ;
		RECT	14.23 411.655 14.28 411.785 ;
		RECT	14.23 413.385 14.28 413.515 ;
		RECT	14.87 413.615 14.92 413.745 ;
		RECT	6.215 413.845 6.265 413.975 ;
		RECT	6.605 413.845 6.655 413.975 ;
		RECT	7.265 413.845 7.315 413.975 ;
		RECT	8.96 413.845 9.01 413.975 ;
		RECT	9.31 413.845 9.36 413.975 ;
		RECT	12.095 413.845 12.145 413.975 ;
		RECT	12.355 413.845 12.405 413.975 ;
		RECT	13.06 413.845 13.11 413.975 ;
		RECT	14.52 413.845 14.57 413.975 ;
		RECT	14.87 229.755 14.92 229.885 ;
		RECT	6.76 230.215 6.81 230.345 ;
		RECT	8.04 230.215 8.09 230.345 ;
		RECT	9.58 230.215 9.63 230.345 ;
		RECT	9.855 230.215 9.905 230.345 ;
		RECT	10.26 230.215 10.31 230.345 ;
		RECT	11.565 230.215 11.615 230.345 ;
		RECT	13.33 230.215 13.38 230.345 ;
		RECT	14.23 230.215 14.28 230.345 ;
		RECT	14.23 231.945 14.28 232.075 ;
		RECT	14.87 232.175 14.92 232.305 ;
		RECT	6.215 232.405 6.265 232.535 ;
		RECT	6.605 232.405 6.655 232.535 ;
		RECT	7.265 232.405 7.315 232.535 ;
		RECT	8.96 232.405 9.01 232.535 ;
		RECT	9.31 232.405 9.36 232.535 ;
		RECT	12.095 232.405 12.145 232.535 ;
		RECT	12.355 232.405 12.405 232.535 ;
		RECT	13.06 232.405 13.11 232.535 ;
		RECT	14.52 232.405 14.57 232.535 ;
		RECT	14.52 414.535 14.57 414.665 ;
		RECT	3.6 414.075 3.65 414.205 ;
		RECT	1.44 414.535 1.49 414.665 ;
		RECT	2.11 414.535 2.16 414.665 ;
		RECT	3.09 414.535 3.14 414.665 ;
		RECT	4.38 414.535 4.43 414.665 ;
		RECT	6.175 414.535 6.225 414.665 ;
		RECT	7.73 414.535 7.78 414.665 ;
		RECT	14.68 414.535 14.73 414.665 ;
		RECT	14.34 414.305 14.39 414.435 ;
		RECT	9.1 414.075 9.15 414.205 ;
		RECT	10.81 414.075 10.86 414.205 ;
		RECT	0.435 414.075 0.485 414.205 ;
		RECT	0.62 414.535 0.67 414.665 ;
		RECT	4.19 414.535 4.24 414.665 ;
		RECT	2.72 414.075 2.77 414.205 ;
		RECT	0.9 235.285 0.95 235.415 ;
		RECT	0.9 261.205 0.95 261.335 ;
		RECT	0.9 264.085 0.95 264.215 ;
		RECT	0.9 266.965 0.95 267.095 ;
		RECT	0.9 269.845 0.95 269.975 ;
		RECT	0.9 272.725 0.95 272.855 ;
		RECT	0.9 275.605 0.95 275.735 ;
		RECT	0.9 278.485 0.95 278.615 ;
		RECT	0.9 281.365 0.95 281.495 ;
		RECT	0.9 284.245 0.95 284.375 ;
		RECT	0.9 287.125 0.95 287.255 ;
		RECT	0.9 238.165 0.95 238.295 ;
		RECT	0.9 290.005 0.95 290.135 ;
		RECT	0.9 292.885 0.95 293.015 ;
		RECT	0.9 295.765 0.95 295.895 ;
		RECT	0.9 298.645 0.95 298.775 ;
		RECT	0.9 301.525 0.95 301.655 ;
		RECT	0.9 304.405 0.95 304.535 ;
		RECT	0.9 307.285 0.95 307.415 ;
		RECT	0.9 310.165 0.95 310.295 ;
		RECT	0.9 313.045 0.95 313.175 ;
		RECT	0.9 315.925 0.95 316.055 ;
		RECT	0.9 241.045 0.95 241.175 ;
		RECT	0.9 318.805 0.95 318.935 ;
		RECT	0.9 321.685 0.95 321.815 ;
		RECT	0.9 324.565 0.95 324.695 ;
		RECT	0.9 327.445 0.95 327.575 ;
		RECT	0.9 330.325 0.95 330.455 ;
		RECT	0.9 333.205 0.95 333.335 ;
		RECT	0.9 336.085 0.95 336.215 ;
		RECT	0.9 338.965 0.95 339.095 ;
		RECT	0.9 341.845 0.95 341.975 ;
		RECT	0.9 344.725 0.95 344.855 ;
		RECT	0.9 243.925 0.95 244.055 ;
		RECT	0.9 347.605 0.95 347.735 ;
		RECT	0.9 350.485 0.95 350.615 ;
		RECT	0.9 353.365 0.95 353.495 ;
		RECT	0.9 356.245 0.95 356.375 ;
		RECT	0.9 359.125 0.95 359.255 ;
		RECT	0.9 362.005 0.95 362.135 ;
		RECT	0.9 364.885 0.95 365.015 ;
		RECT	0.9 367.765 0.95 367.895 ;
		RECT	0.9 370.645 0.95 370.775 ;
		RECT	0.9 373.525 0.95 373.655 ;
		RECT	0.9 246.805 0.95 246.935 ;
		RECT	0.9 376.405 0.95 376.535 ;
		RECT	0.9 379.285 0.95 379.415 ;
		RECT	0.9 382.165 0.95 382.295 ;
		RECT	0.9 385.045 0.95 385.175 ;
		RECT	0.9 387.925 0.95 388.055 ;
		RECT	0.9 390.805 0.95 390.935 ;
		RECT	0.9 393.685 0.95 393.815 ;
		RECT	0.9 396.565 0.95 396.695 ;
		RECT	0.9 399.445 0.95 399.575 ;
		RECT	0.9 402.325 0.95 402.455 ;
		RECT	0.9 249.685 0.95 249.815 ;
		RECT	0.9 405.205 0.95 405.335 ;
		RECT	0.9 408.085 0.95 408.215 ;
		RECT	0.9 410.965 0.95 411.095 ;
		RECT	0.9 252.565 0.95 252.695 ;
		RECT	0.9 255.445 0.95 255.575 ;
		RECT	0.9 258.325 0.95 258.455 ;
		RECT	0.9 413.845 0.95 413.975 ;
		RECT	0.9 232.405 0.95 232.535 ;
		RECT	2.72 229.755 2.77 229.885 ;
		RECT	2.72 232.175 2.77 232.305 ;
		RECT	2.72 258.555 2.77 258.685 ;
		RECT	2.72 260.975 2.77 261.105 ;
		RECT	2.72 261.435 2.77 261.565 ;
		RECT	2.72 263.855 2.77 263.985 ;
		RECT	2.72 264.315 2.77 264.445 ;
		RECT	2.72 266.735 2.77 266.865 ;
		RECT	2.72 267.195 2.77 267.325 ;
		RECT	2.72 269.615 2.77 269.745 ;
		RECT	2.72 270.075 2.77 270.205 ;
		RECT	2.72 272.495 2.77 272.625 ;
		RECT	2.72 272.955 2.77 273.085 ;
		RECT	2.72 275.375 2.77 275.505 ;
		RECT	2.72 275.835 2.77 275.965 ;
		RECT	2.72 278.255 2.77 278.385 ;
		RECT	2.72 278.715 2.77 278.845 ;
		RECT	2.72 281.135 2.77 281.265 ;
		RECT	2.72 281.595 2.77 281.725 ;
		RECT	2.72 284.015 2.77 284.145 ;
		RECT	2.72 284.475 2.77 284.605 ;
		RECT	2.72 286.895 2.77 287.025 ;
		RECT	2.72 232.635 2.77 232.765 ;
		RECT	2.72 235.055 2.77 235.185 ;
		RECT	2.72 287.355 2.77 287.485 ;
		RECT	2.72 289.775 2.77 289.905 ;
		RECT	2.72 290.235 2.77 290.365 ;
		RECT	2.72 292.655 2.77 292.785 ;
		RECT	2.72 293.115 2.77 293.245 ;
		RECT	2.72 295.535 2.77 295.665 ;
		RECT	2.72 295.995 2.77 296.125 ;
		RECT	2.72 298.415 2.77 298.545 ;
		RECT	2.72 298.875 2.77 299.005 ;
		RECT	2.72 301.295 2.77 301.425 ;
		RECT	2.72 301.755 2.77 301.885 ;
		RECT	2.72 304.175 2.77 304.305 ;
		RECT	2.72 304.635 2.77 304.765 ;
		RECT	2.72 307.055 2.77 307.185 ;
		RECT	2.72 307.515 2.77 307.645 ;
		RECT	2.72 309.935 2.77 310.065 ;
		RECT	2.72 310.395 2.77 310.525 ;
		RECT	2.72 312.815 2.77 312.945 ;
		RECT	2.72 313.275 2.77 313.405 ;
		RECT	2.72 315.695 2.77 315.825 ;
		RECT	2.72 235.515 2.77 235.645 ;
		RECT	2.72 237.935 2.77 238.065 ;
		RECT	2.72 316.155 2.77 316.285 ;
		RECT	2.72 318.575 2.77 318.705 ;
		RECT	2.72 319.035 2.77 319.165 ;
		RECT	2.72 321.455 2.77 321.585 ;
		RECT	2.72 321.915 2.77 322.045 ;
		RECT	2.72 324.335 2.77 324.465 ;
		RECT	2.72 324.795 2.77 324.925 ;
		RECT	2.72 327.215 2.77 327.345 ;
		RECT	2.72 327.675 2.77 327.805 ;
		RECT	2.72 330.095 2.77 330.225 ;
		RECT	2.72 330.555 2.77 330.685 ;
		RECT	2.72 332.975 2.77 333.105 ;
		RECT	2.72 333.435 2.77 333.565 ;
		RECT	2.72 335.855 2.77 335.985 ;
		RECT	2.72 336.315 2.77 336.445 ;
		RECT	2.72 338.735 2.77 338.865 ;
		RECT	2.72 339.195 2.77 339.325 ;
		RECT	2.72 341.615 2.77 341.745 ;
		RECT	2.72 342.075 2.77 342.205 ;
		RECT	2.72 344.495 2.77 344.625 ;
		RECT	2.72 238.395 2.77 238.525 ;
		RECT	2.72 240.815 2.77 240.945 ;
		RECT	2.72 344.955 2.77 345.085 ;
		RECT	2.72 347.375 2.77 347.505 ;
		RECT	2.72 347.835 2.77 347.965 ;
		RECT	2.72 350.255 2.77 350.385 ;
		RECT	2.72 350.715 2.77 350.845 ;
		RECT	2.72 353.135 2.77 353.265 ;
		RECT	2.72 353.595 2.77 353.725 ;
		RECT	2.72 356.015 2.77 356.145 ;
		RECT	2.72 356.475 2.77 356.605 ;
		RECT	2.72 358.895 2.77 359.025 ;
		RECT	2.72 359.355 2.77 359.485 ;
		RECT	2.72 361.775 2.77 361.905 ;
		RECT	2.72 362.235 2.77 362.365 ;
		RECT	2.72 364.655 2.77 364.785 ;
		RECT	2.72 365.115 2.77 365.245 ;
		RECT	2.72 367.535 2.77 367.665 ;
		RECT	2.72 367.995 2.77 368.125 ;
		RECT	2.72 370.415 2.77 370.545 ;
		RECT	2.72 370.875 2.77 371.005 ;
		RECT	2.72 373.295 2.77 373.425 ;
		RECT	2.72 241.275 2.77 241.405 ;
		RECT	2.72 243.695 2.77 243.825 ;
		RECT	2.72 373.755 2.77 373.885 ;
		RECT	2.72 376.175 2.77 376.305 ;
		RECT	2.72 376.635 2.77 376.765 ;
		RECT	2.72 379.055 2.77 379.185 ;
		RECT	2.72 379.515 2.77 379.645 ;
		RECT	2.72 381.935 2.77 382.065 ;
		RECT	2.72 382.395 2.77 382.525 ;
		RECT	2.72 384.815 2.77 384.945 ;
		RECT	2.72 385.275 2.77 385.405 ;
		RECT	2.72 387.695 2.77 387.825 ;
		RECT	2.72 388.155 2.77 388.285 ;
		RECT	2.72 390.575 2.77 390.705 ;
		RECT	2.72 391.035 2.77 391.165 ;
		RECT	2.72 393.455 2.77 393.585 ;
		RECT	2.72 393.915 2.77 394.045 ;
		RECT	2.72 396.335 2.77 396.465 ;
		RECT	2.72 396.795 2.77 396.925 ;
		RECT	2.72 399.215 2.77 399.345 ;
		RECT	2.72 399.675 2.77 399.805 ;
		RECT	2.72 402.095 2.77 402.225 ;
		RECT	2.72 244.155 2.77 244.285 ;
		RECT	2.72 246.575 2.77 246.705 ;
		RECT	2.72 402.555 2.77 402.685 ;
		RECT	2.72 404.975 2.77 405.105 ;
		RECT	2.72 405.435 2.77 405.565 ;
		RECT	2.72 407.855 2.77 407.985 ;
		RECT	2.72 408.315 2.77 408.445 ;
		RECT	2.72 410.735 2.77 410.865 ;
		RECT	2.72 411.195 2.77 411.325 ;
		RECT	2.72 413.615 2.77 413.745 ;
		RECT	2.72 247.035 2.77 247.165 ;
		RECT	2.72 249.455 2.77 249.585 ;
		RECT	2.72 249.915 2.77 250.045 ;
		RECT	2.72 252.335 2.77 252.465 ;
		RECT	2.72 252.795 2.77 252.925 ;
		RECT	2.72 255.215 2.77 255.345 ;
		RECT	2.72 255.675 2.77 255.805 ;
		RECT	2.72 258.095 2.77 258.225 ;
		RECT	1.625 229.755 1.675 229.885 ;
		RECT	1.92 229.755 1.97 229.885 ;
		RECT	5.05 229.755 5.1 229.885 ;
		RECT	3.6 230.215 3.65 230.345 ;
		RECT	1.625 232.175 1.675 232.305 ;
		RECT	1.92 232.175 1.97 232.305 ;
		RECT	5.05 232.175 5.1 232.305 ;
		RECT	1.625 258.555 1.675 258.685 ;
		RECT	1.92 258.555 1.97 258.685 ;
		RECT	5.05 258.555 5.1 258.685 ;
		RECT	3.6 259.015 3.65 259.145 ;
		RECT	1.625 260.975 1.675 261.105 ;
		RECT	1.92 260.975 1.97 261.105 ;
		RECT	5.05 260.975 5.1 261.105 ;
		RECT	1.625 261.435 1.675 261.565 ;
		RECT	1.92 261.435 1.97 261.565 ;
		RECT	5.05 261.435 5.1 261.565 ;
		RECT	3.6 261.895 3.65 262.025 ;
		RECT	1.625 263.855 1.675 263.985 ;
		RECT	1.92 263.855 1.97 263.985 ;
		RECT	5.05 263.855 5.1 263.985 ;
		RECT	1.625 264.315 1.675 264.445 ;
		RECT	1.92 264.315 1.97 264.445 ;
		RECT	5.05 264.315 5.1 264.445 ;
		RECT	3.6 264.775 3.65 264.905 ;
		RECT	1.625 266.735 1.675 266.865 ;
		RECT	1.92 266.735 1.97 266.865 ;
		RECT	5.05 266.735 5.1 266.865 ;
		RECT	1.625 267.195 1.675 267.325 ;
		RECT	1.92 267.195 1.97 267.325 ;
		RECT	5.05 267.195 5.1 267.325 ;
		RECT	3.6 267.655 3.65 267.785 ;
		RECT	1.625 269.615 1.675 269.745 ;
		RECT	1.92 269.615 1.97 269.745 ;
		RECT	5.05 269.615 5.1 269.745 ;
		RECT	1.625 270.075 1.675 270.205 ;
		RECT	1.92 270.075 1.97 270.205 ;
		RECT	5.05 270.075 5.1 270.205 ;
		RECT	3.6 270.535 3.65 270.665 ;
		RECT	1.625 272.495 1.675 272.625 ;
		RECT	1.92 272.495 1.97 272.625 ;
		RECT	5.05 272.495 5.1 272.625 ;
		RECT	1.625 272.955 1.675 273.085 ;
		RECT	1.92 272.955 1.97 273.085 ;
		RECT	5.05 272.955 5.1 273.085 ;
		RECT	3.6 273.415 3.65 273.545 ;
		RECT	1.625 275.375 1.675 275.505 ;
		RECT	1.92 275.375 1.97 275.505 ;
		RECT	5.05 275.375 5.1 275.505 ;
		RECT	1.625 275.835 1.675 275.965 ;
		RECT	1.92 275.835 1.97 275.965 ;
		RECT	5.05 275.835 5.1 275.965 ;
		RECT	3.6 276.295 3.65 276.425 ;
		RECT	1.625 278.255 1.675 278.385 ;
		RECT	1.92 278.255 1.97 278.385 ;
		RECT	5.05 278.255 5.1 278.385 ;
		RECT	1.625 278.715 1.675 278.845 ;
		RECT	1.92 278.715 1.97 278.845 ;
		RECT	5.05 278.715 5.1 278.845 ;
		RECT	3.6 279.175 3.65 279.305 ;
		RECT	1.625 281.135 1.675 281.265 ;
		RECT	1.92 281.135 1.97 281.265 ;
		RECT	5.05 281.135 5.1 281.265 ;
		RECT	1.625 281.595 1.675 281.725 ;
		RECT	1.92 281.595 1.97 281.725 ;
		RECT	5.05 281.595 5.1 281.725 ;
		RECT	3.6 282.055 3.65 282.185 ;
		RECT	1.625 284.015 1.675 284.145 ;
		RECT	1.92 284.015 1.97 284.145 ;
		RECT	5.05 284.015 5.1 284.145 ;
		RECT	1.625 284.475 1.675 284.605 ;
		RECT	1.92 284.475 1.97 284.605 ;
		RECT	5.05 284.475 5.1 284.605 ;
		RECT	3.6 284.935 3.65 285.065 ;
		RECT	1.625 286.895 1.675 287.025 ;
		RECT	1.92 286.895 1.97 287.025 ;
		RECT	5.05 286.895 5.1 287.025 ;
		RECT	1.625 232.635 1.675 232.765 ;
		RECT	1.92 232.635 1.97 232.765 ;
		RECT	5.05 232.635 5.1 232.765 ;
		RECT	3.6 233.095 3.65 233.225 ;
		RECT	1.625 235.055 1.675 235.185 ;
		RECT	1.92 235.055 1.97 235.185 ;
		RECT	5.05 235.055 5.1 235.185 ;
		RECT	1.625 287.355 1.675 287.485 ;
		RECT	1.92 287.355 1.97 287.485 ;
		RECT	5.05 287.355 5.1 287.485 ;
		RECT	3.6 287.815 3.65 287.945 ;
		RECT	1.625 289.775 1.675 289.905 ;
		RECT	1.92 289.775 1.97 289.905 ;
		RECT	5.05 289.775 5.1 289.905 ;
		RECT	1.625 290.235 1.675 290.365 ;
		RECT	1.92 290.235 1.97 290.365 ;
		RECT	5.05 290.235 5.1 290.365 ;
		RECT	3.6 290.695 3.65 290.825 ;
		RECT	1.625 292.655 1.675 292.785 ;
		RECT	1.92 292.655 1.97 292.785 ;
		RECT	5.05 292.655 5.1 292.785 ;
		RECT	1.625 293.115 1.675 293.245 ;
		RECT	1.92 293.115 1.97 293.245 ;
		RECT	5.05 293.115 5.1 293.245 ;
		RECT	3.6 293.575 3.65 293.705 ;
		RECT	1.625 295.535 1.675 295.665 ;
		RECT	1.92 295.535 1.97 295.665 ;
		RECT	5.05 295.535 5.1 295.665 ;
		RECT	1.625 295.995 1.675 296.125 ;
		RECT	1.92 295.995 1.97 296.125 ;
		RECT	5.05 295.995 5.1 296.125 ;
		RECT	3.6 296.455 3.65 296.585 ;
		RECT	1.625 298.415 1.675 298.545 ;
		RECT	1.92 298.415 1.97 298.545 ;
		RECT	5.05 298.415 5.1 298.545 ;
		RECT	1.625 298.875 1.675 299.005 ;
		RECT	1.92 298.875 1.97 299.005 ;
		RECT	5.05 298.875 5.1 299.005 ;
		RECT	3.6 299.335 3.65 299.465 ;
		RECT	1.625 301.295 1.675 301.425 ;
		RECT	1.92 301.295 1.97 301.425 ;
		RECT	5.05 301.295 5.1 301.425 ;
		RECT	1.625 301.755 1.675 301.885 ;
		RECT	1.92 301.755 1.97 301.885 ;
		RECT	5.05 301.755 5.1 301.885 ;
		RECT	3.6 302.215 3.65 302.345 ;
		RECT	1.625 304.175 1.675 304.305 ;
		RECT	1.92 304.175 1.97 304.305 ;
		RECT	5.05 304.175 5.1 304.305 ;
		RECT	1.625 304.635 1.675 304.765 ;
		RECT	1.92 304.635 1.97 304.765 ;
		RECT	5.05 304.635 5.1 304.765 ;
		RECT	3.6 305.095 3.65 305.225 ;
		RECT	1.625 307.055 1.675 307.185 ;
		RECT	1.92 307.055 1.97 307.185 ;
		RECT	5.05 307.055 5.1 307.185 ;
		RECT	1.625 307.515 1.675 307.645 ;
		RECT	1.92 307.515 1.97 307.645 ;
		RECT	5.05 307.515 5.1 307.645 ;
		RECT	3.6 307.975 3.65 308.105 ;
		RECT	1.625 309.935 1.675 310.065 ;
		RECT	1.92 309.935 1.97 310.065 ;
		RECT	5.05 309.935 5.1 310.065 ;
		RECT	1.625 310.395 1.675 310.525 ;
		RECT	1.92 310.395 1.97 310.525 ;
		RECT	5.05 310.395 5.1 310.525 ;
		RECT	3.6 310.855 3.65 310.985 ;
		RECT	1.625 312.815 1.675 312.945 ;
		RECT	1.92 312.815 1.97 312.945 ;
		RECT	5.05 312.815 5.1 312.945 ;
		RECT	1.625 313.275 1.675 313.405 ;
		RECT	1.92 313.275 1.97 313.405 ;
		RECT	5.05 313.275 5.1 313.405 ;
		RECT	3.6 313.735 3.65 313.865 ;
		RECT	1.625 315.695 1.675 315.825 ;
		RECT	1.92 315.695 1.97 315.825 ;
		RECT	5.05 315.695 5.1 315.825 ;
		RECT	1.625 235.515 1.675 235.645 ;
		RECT	1.92 235.515 1.97 235.645 ;
		RECT	5.05 235.515 5.1 235.645 ;
		RECT	3.6 235.975 3.65 236.105 ;
		RECT	1.625 237.935 1.675 238.065 ;
		RECT	1.92 237.935 1.97 238.065 ;
		RECT	5.05 237.935 5.1 238.065 ;
		RECT	1.625 316.155 1.675 316.285 ;
		RECT	1.92 316.155 1.97 316.285 ;
		RECT	5.05 316.155 5.1 316.285 ;
		RECT	3.6 316.615 3.65 316.745 ;
		RECT	1.625 318.575 1.675 318.705 ;
		RECT	1.92 318.575 1.97 318.705 ;
		RECT	5.05 318.575 5.1 318.705 ;
		RECT	1.625 319.035 1.675 319.165 ;
		RECT	1.92 319.035 1.97 319.165 ;
		RECT	5.05 319.035 5.1 319.165 ;
		RECT	3.6 319.495 3.65 319.625 ;
		RECT	1.625 321.455 1.675 321.585 ;
		RECT	1.92 321.455 1.97 321.585 ;
		RECT	5.05 321.455 5.1 321.585 ;
		RECT	1.625 321.915 1.675 322.045 ;
		RECT	1.92 321.915 1.97 322.045 ;
		RECT	5.05 321.915 5.1 322.045 ;
		RECT	3.6 322.375 3.65 322.505 ;
		RECT	1.625 324.335 1.675 324.465 ;
		RECT	1.92 324.335 1.97 324.465 ;
		RECT	5.05 324.335 5.1 324.465 ;
		RECT	1.625 324.795 1.675 324.925 ;
		RECT	1.92 324.795 1.97 324.925 ;
		RECT	5.05 324.795 5.1 324.925 ;
		RECT	3.6 325.255 3.65 325.385 ;
		RECT	1.625 327.215 1.675 327.345 ;
		RECT	1.92 327.215 1.97 327.345 ;
		RECT	5.05 327.215 5.1 327.345 ;
		RECT	1.625 327.675 1.675 327.805 ;
		RECT	1.92 327.675 1.97 327.805 ;
		RECT	5.05 327.675 5.1 327.805 ;
		RECT	3.6 328.135 3.65 328.265 ;
		RECT	1.625 330.095 1.675 330.225 ;
		RECT	1.92 330.095 1.97 330.225 ;
		RECT	5.05 330.095 5.1 330.225 ;
		RECT	1.625 330.555 1.675 330.685 ;
		RECT	1.92 330.555 1.97 330.685 ;
		RECT	5.05 330.555 5.1 330.685 ;
		RECT	3.6 331.015 3.65 331.145 ;
		RECT	1.625 332.975 1.675 333.105 ;
		RECT	1.92 332.975 1.97 333.105 ;
		RECT	5.05 332.975 5.1 333.105 ;
		RECT	1.625 333.435 1.675 333.565 ;
		RECT	1.92 333.435 1.97 333.565 ;
		RECT	5.05 333.435 5.1 333.565 ;
		RECT	3.6 333.895 3.65 334.025 ;
		RECT	1.625 335.855 1.675 335.985 ;
		RECT	1.92 335.855 1.97 335.985 ;
		RECT	5.05 335.855 5.1 335.985 ;
		RECT	1.625 336.315 1.675 336.445 ;
		RECT	1.92 336.315 1.97 336.445 ;
		RECT	5.05 336.315 5.1 336.445 ;
		RECT	3.6 336.775 3.65 336.905 ;
		RECT	1.625 338.735 1.675 338.865 ;
		RECT	1.92 338.735 1.97 338.865 ;
		RECT	5.05 338.735 5.1 338.865 ;
		RECT	1.625 339.195 1.675 339.325 ;
		RECT	1.92 339.195 1.97 339.325 ;
		RECT	5.05 339.195 5.1 339.325 ;
		RECT	3.6 339.655 3.65 339.785 ;
		RECT	1.625 341.615 1.675 341.745 ;
		RECT	1.92 341.615 1.97 341.745 ;
		RECT	5.05 341.615 5.1 341.745 ;
		RECT	1.625 342.075 1.675 342.205 ;
		RECT	1.92 342.075 1.97 342.205 ;
		RECT	5.05 342.075 5.1 342.205 ;
		RECT	3.6 342.535 3.65 342.665 ;
		RECT	1.625 344.495 1.675 344.625 ;
		RECT	1.92 344.495 1.97 344.625 ;
		RECT	5.05 344.495 5.1 344.625 ;
		RECT	1.625 238.395 1.675 238.525 ;
		RECT	1.92 238.395 1.97 238.525 ;
		RECT	5.05 238.395 5.1 238.525 ;
		RECT	3.6 238.855 3.65 238.985 ;
		RECT	1.625 240.815 1.675 240.945 ;
		RECT	1.92 240.815 1.97 240.945 ;
		RECT	5.05 240.815 5.1 240.945 ;
		RECT	1.625 344.955 1.675 345.085 ;
		RECT	1.92 344.955 1.97 345.085 ;
		RECT	5.05 344.955 5.1 345.085 ;
		RECT	3.6 345.415 3.65 345.545 ;
		RECT	1.625 347.375 1.675 347.505 ;
		RECT	1.92 347.375 1.97 347.505 ;
		RECT	5.05 347.375 5.1 347.505 ;
		RECT	1.625 347.835 1.675 347.965 ;
		RECT	1.92 347.835 1.97 347.965 ;
		RECT	5.05 347.835 5.1 347.965 ;
		RECT	3.6 348.295 3.65 348.425 ;
		RECT	1.625 350.255 1.675 350.385 ;
		RECT	1.92 350.255 1.97 350.385 ;
		RECT	5.05 350.255 5.1 350.385 ;
		RECT	1.625 350.715 1.675 350.845 ;
		RECT	1.92 350.715 1.97 350.845 ;
		RECT	5.05 350.715 5.1 350.845 ;
		RECT	3.6 351.175 3.65 351.305 ;
		RECT	1.625 353.135 1.675 353.265 ;
		RECT	1.92 353.135 1.97 353.265 ;
		RECT	5.05 353.135 5.1 353.265 ;
		RECT	1.625 353.595 1.675 353.725 ;
		RECT	1.92 353.595 1.97 353.725 ;
		RECT	5.05 353.595 5.1 353.725 ;
		RECT	3.6 354.055 3.65 354.185 ;
		RECT	1.625 356.015 1.675 356.145 ;
		RECT	1.92 356.015 1.97 356.145 ;
		RECT	5.05 356.015 5.1 356.145 ;
		RECT	1.625 356.475 1.675 356.605 ;
		RECT	1.92 356.475 1.97 356.605 ;
		RECT	5.05 356.475 5.1 356.605 ;
		RECT	3.6 356.935 3.65 357.065 ;
		RECT	1.625 358.895 1.675 359.025 ;
		RECT	1.92 358.895 1.97 359.025 ;
		RECT	5.05 358.895 5.1 359.025 ;
		RECT	1.625 359.355 1.675 359.485 ;
		RECT	1.92 359.355 1.97 359.485 ;
		RECT	5.05 359.355 5.1 359.485 ;
		RECT	3.6 359.815 3.65 359.945 ;
		RECT	1.625 361.775 1.675 361.905 ;
		RECT	1.92 361.775 1.97 361.905 ;
		RECT	5.05 361.775 5.1 361.905 ;
		RECT	1.625 362.235 1.675 362.365 ;
		RECT	1.92 362.235 1.97 362.365 ;
		RECT	5.05 362.235 5.1 362.365 ;
		RECT	3.6 362.695 3.65 362.825 ;
		RECT	1.625 364.655 1.675 364.785 ;
		RECT	1.92 364.655 1.97 364.785 ;
		RECT	5.05 364.655 5.1 364.785 ;
		RECT	1.625 365.115 1.675 365.245 ;
		RECT	1.92 365.115 1.97 365.245 ;
		RECT	5.05 365.115 5.1 365.245 ;
		RECT	3.6 365.575 3.65 365.705 ;
		RECT	1.625 367.535 1.675 367.665 ;
		RECT	1.92 367.535 1.97 367.665 ;
		RECT	5.05 367.535 5.1 367.665 ;
		RECT	1.625 367.995 1.675 368.125 ;
		RECT	1.92 367.995 1.97 368.125 ;
		RECT	5.05 367.995 5.1 368.125 ;
		RECT	3.6 368.455 3.65 368.585 ;
		RECT	1.625 370.415 1.675 370.545 ;
		RECT	1.92 370.415 1.97 370.545 ;
		RECT	5.05 370.415 5.1 370.545 ;
		RECT	1.625 370.875 1.675 371.005 ;
		RECT	1.92 370.875 1.97 371.005 ;
		RECT	5.05 370.875 5.1 371.005 ;
		RECT	3.6 371.335 3.65 371.465 ;
		RECT	1.625 373.295 1.675 373.425 ;
		RECT	1.92 373.295 1.97 373.425 ;
		RECT	5.05 373.295 5.1 373.425 ;
		RECT	1.625 241.275 1.675 241.405 ;
		RECT	1.92 241.275 1.97 241.405 ;
		RECT	5.05 241.275 5.1 241.405 ;
		RECT	3.6 241.735 3.65 241.865 ;
		RECT	1.625 243.695 1.675 243.825 ;
		RECT	1.92 243.695 1.97 243.825 ;
		RECT	5.05 243.695 5.1 243.825 ;
		RECT	1.625 373.755 1.675 373.885 ;
		RECT	1.92 373.755 1.97 373.885 ;
		RECT	5.05 373.755 5.1 373.885 ;
		RECT	3.6 374.215 3.65 374.345 ;
		RECT	1.625 376.175 1.675 376.305 ;
		RECT	1.92 376.175 1.97 376.305 ;
		RECT	5.05 376.175 5.1 376.305 ;
		RECT	1.625 376.635 1.675 376.765 ;
		RECT	1.92 376.635 1.97 376.765 ;
		RECT	5.05 376.635 5.1 376.765 ;
		RECT	3.6 377.095 3.65 377.225 ;
		RECT	1.625 379.055 1.675 379.185 ;
		RECT	1.92 379.055 1.97 379.185 ;
		RECT	5.05 379.055 5.1 379.185 ;
		RECT	1.625 379.515 1.675 379.645 ;
		RECT	1.92 379.515 1.97 379.645 ;
		RECT	5.05 379.515 5.1 379.645 ;
		RECT	3.6 379.975 3.65 380.105 ;
		RECT	1.625 381.935 1.675 382.065 ;
		RECT	1.92 381.935 1.97 382.065 ;
		RECT	5.05 381.935 5.1 382.065 ;
		RECT	1.625 382.395 1.675 382.525 ;
		RECT	1.92 382.395 1.97 382.525 ;
		RECT	5.05 382.395 5.1 382.525 ;
		RECT	3.6 382.855 3.65 382.985 ;
		RECT	1.625 384.815 1.675 384.945 ;
		RECT	1.92 384.815 1.97 384.945 ;
		RECT	5.05 384.815 5.1 384.945 ;
		RECT	1.625 385.275 1.675 385.405 ;
		RECT	1.92 385.275 1.97 385.405 ;
		RECT	5.05 385.275 5.1 385.405 ;
		RECT	3.6 385.735 3.65 385.865 ;
		RECT	1.625 387.695 1.675 387.825 ;
		RECT	1.92 387.695 1.97 387.825 ;
		RECT	5.05 387.695 5.1 387.825 ;
		RECT	1.625 388.155 1.675 388.285 ;
		RECT	1.92 388.155 1.97 388.285 ;
		RECT	5.05 388.155 5.1 388.285 ;
		RECT	3.6 388.615 3.65 388.745 ;
		RECT	1.625 390.575 1.675 390.705 ;
		RECT	1.92 390.575 1.97 390.705 ;
		RECT	5.05 390.575 5.1 390.705 ;
		RECT	1.625 391.035 1.675 391.165 ;
		RECT	1.92 391.035 1.97 391.165 ;
		RECT	5.05 391.035 5.1 391.165 ;
		RECT	3.6 391.495 3.65 391.625 ;
		RECT	1.625 393.455 1.675 393.585 ;
		RECT	1.92 393.455 1.97 393.585 ;
		RECT	5.05 393.455 5.1 393.585 ;
		RECT	1.625 393.915 1.675 394.045 ;
		RECT	1.92 393.915 1.97 394.045 ;
		RECT	5.05 393.915 5.1 394.045 ;
		RECT	3.6 394.375 3.65 394.505 ;
		RECT	1.625 396.335 1.675 396.465 ;
		RECT	1.92 396.335 1.97 396.465 ;
		RECT	5.05 396.335 5.1 396.465 ;
		RECT	1.625 396.795 1.675 396.925 ;
		RECT	1.92 396.795 1.97 396.925 ;
		RECT	5.05 396.795 5.1 396.925 ;
		RECT	3.6 397.255 3.65 397.385 ;
		RECT	1.625 399.215 1.675 399.345 ;
		RECT	1.92 399.215 1.97 399.345 ;
		RECT	5.05 399.215 5.1 399.345 ;
		RECT	1.625 399.675 1.675 399.805 ;
		RECT	1.92 399.675 1.97 399.805 ;
		RECT	5.05 399.675 5.1 399.805 ;
		RECT	3.6 400.135 3.65 400.265 ;
		RECT	1.625 402.095 1.675 402.225 ;
		RECT	1.92 402.095 1.97 402.225 ;
		RECT	5.05 402.095 5.1 402.225 ;
		RECT	1.625 244.155 1.675 244.285 ;
		RECT	1.92 244.155 1.97 244.285 ;
		RECT	5.05 244.155 5.1 244.285 ;
		RECT	3.6 244.615 3.65 244.745 ;
		RECT	1.625 246.575 1.675 246.705 ;
		RECT	1.92 246.575 1.97 246.705 ;
		RECT	5.05 246.575 5.1 246.705 ;
		RECT	1.625 402.555 1.675 402.685 ;
		RECT	1.92 402.555 1.97 402.685 ;
		RECT	5.05 402.555 5.1 402.685 ;
		RECT	3.6 403.015 3.65 403.145 ;
		RECT	1.625 404.975 1.675 405.105 ;
		RECT	1.92 404.975 1.97 405.105 ;
		RECT	5.05 404.975 5.1 405.105 ;
		RECT	1.625 405.435 1.675 405.565 ;
		RECT	1.92 405.435 1.97 405.565 ;
		RECT	5.05 405.435 5.1 405.565 ;
		RECT	3.6 405.895 3.65 406.025 ;
		RECT	1.625 407.855 1.675 407.985 ;
		RECT	1.92 407.855 1.97 407.985 ;
		RECT	5.05 407.855 5.1 407.985 ;
		RECT	1.625 408.315 1.675 408.445 ;
		RECT	1.92 408.315 1.97 408.445 ;
		RECT	5.05 408.315 5.1 408.445 ;
		RECT	3.6 408.775 3.65 408.905 ;
		RECT	1.625 410.735 1.675 410.865 ;
		RECT	1.92 410.735 1.97 410.865 ;
		RECT	5.05 410.735 5.1 410.865 ;
		RECT	1.625 411.195 1.675 411.325 ;
		RECT	1.92 411.195 1.97 411.325 ;
		RECT	5.05 411.195 5.1 411.325 ;
		RECT	3.6 411.655 3.65 411.785 ;
		RECT	1.625 413.615 1.675 413.745 ;
		RECT	1.92 413.615 1.97 413.745 ;
		RECT	5.05 413.615 5.1 413.745 ;
		RECT	1.625 247.035 1.675 247.165 ;
		RECT	1.92 247.035 1.97 247.165 ;
		RECT	5.05 247.035 5.1 247.165 ;
		RECT	3.6 247.495 3.65 247.625 ;
		RECT	1.625 249.455 1.675 249.585 ;
		RECT	1.92 249.455 1.97 249.585 ;
		RECT	5.05 249.455 5.1 249.585 ;
		RECT	1.625 249.915 1.675 250.045 ;
		RECT	1.92 249.915 1.97 250.045 ;
		RECT	5.05 249.915 5.1 250.045 ;
		RECT	3.6 250.375 3.65 250.505 ;
		RECT	1.625 252.335 1.675 252.465 ;
		RECT	1.92 252.335 1.97 252.465 ;
		RECT	5.05 252.335 5.1 252.465 ;
		RECT	1.625 252.795 1.675 252.925 ;
		RECT	1.92 252.795 1.97 252.925 ;
		RECT	5.05 252.795 5.1 252.925 ;
		RECT	3.6 253.255 3.65 253.385 ;
		RECT	1.625 255.215 1.675 255.345 ;
		RECT	1.92 255.215 1.97 255.345 ;
		RECT	5.05 255.215 5.1 255.345 ;
		RECT	1.625 255.675 1.675 255.805 ;
		RECT	1.92 255.675 1.97 255.805 ;
		RECT	5.05 255.675 5.1 255.805 ;
		RECT	3.6 256.135 3.65 256.265 ;
		RECT	1.625 258.095 1.675 258.225 ;
		RECT	1.92 258.095 1.97 258.225 ;
		RECT	5.05 258.095 5.1 258.225 ;
		RECT	3.6 232.635 3.65 232.765 ;
		RECT	1.625 233.095 1.675 233.225 ;
		RECT	1.88 233.135 2.01 233.185 ;
		RECT	5.01 233.135 5.14 233.185 ;
		RECT	3.6 235.055 3.65 235.185 ;
		RECT	1.44 235.285 1.49 235.415 ;
		RECT	2.11 235.285 2.16 235.415 ;
		RECT	3.09 235.285 3.14 235.415 ;
		RECT	4.38 235.285 4.43 235.415 ;
		RECT	6.215 235.285 6.265 235.415 ;
		RECT	3.6 258.555 3.65 258.685 ;
		RECT	1.625 259.015 1.675 259.145 ;
		RECT	1.88 259.055 2.01 259.105 ;
		RECT	5.01 259.055 5.14 259.105 ;
		RECT	3.6 260.975 3.65 261.105 ;
		RECT	1.44 261.205 1.49 261.335 ;
		RECT	2.11 261.205 2.16 261.335 ;
		RECT	3.09 261.205 3.14 261.335 ;
		RECT	4.38 261.205 4.43 261.335 ;
		RECT	6.215 261.205 6.265 261.335 ;
		RECT	3.6 261.435 3.65 261.565 ;
		RECT	1.625 261.895 1.675 262.025 ;
		RECT	1.88 261.935 2.01 261.985 ;
		RECT	5.01 261.935 5.14 261.985 ;
		RECT	3.6 263.855 3.65 263.985 ;
		RECT	1.44 264.085 1.49 264.215 ;
		RECT	2.11 264.085 2.16 264.215 ;
		RECT	3.09 264.085 3.14 264.215 ;
		RECT	4.38 264.085 4.43 264.215 ;
		RECT	6.215 264.085 6.265 264.215 ;
		RECT	3.6 264.315 3.65 264.445 ;
		RECT	1.625 264.775 1.675 264.905 ;
		RECT	1.88 264.815 2.01 264.865 ;
		RECT	5.01 264.815 5.14 264.865 ;
		RECT	3.6 266.735 3.65 266.865 ;
		RECT	1.44 266.965 1.49 267.095 ;
		RECT	2.11 266.965 2.16 267.095 ;
		RECT	3.09 266.965 3.14 267.095 ;
		RECT	4.38 266.965 4.43 267.095 ;
		RECT	6.215 266.965 6.265 267.095 ;
		RECT	3.6 267.195 3.65 267.325 ;
		RECT	1.625 267.655 1.675 267.785 ;
		RECT	1.88 267.695 2.01 267.745 ;
		RECT	5.01 267.695 5.14 267.745 ;
		RECT	3.6 269.615 3.65 269.745 ;
		RECT	1.44 269.845 1.49 269.975 ;
		RECT	2.11 269.845 2.16 269.975 ;
		RECT	3.09 269.845 3.14 269.975 ;
		RECT	4.38 269.845 4.43 269.975 ;
		RECT	6.215 269.845 6.265 269.975 ;
		RECT	3.6 270.075 3.65 270.205 ;
		RECT	1.625 270.535 1.675 270.665 ;
		RECT	1.88 270.575 2.01 270.625 ;
		RECT	5.01 270.575 5.14 270.625 ;
		RECT	3.6 272.495 3.65 272.625 ;
		RECT	1.44 272.725 1.49 272.855 ;
		RECT	2.11 272.725 2.16 272.855 ;
		RECT	3.09 272.725 3.14 272.855 ;
		RECT	4.38 272.725 4.43 272.855 ;
		RECT	6.215 272.725 6.265 272.855 ;
		RECT	3.6 272.955 3.65 273.085 ;
		RECT	1.625 273.415 1.675 273.545 ;
		RECT	1.88 273.455 2.01 273.505 ;
		RECT	5.01 273.455 5.14 273.505 ;
		RECT	3.6 275.375 3.65 275.505 ;
		RECT	1.44 275.605 1.49 275.735 ;
		RECT	2.11 275.605 2.16 275.735 ;
		RECT	3.09 275.605 3.14 275.735 ;
		RECT	4.38 275.605 4.43 275.735 ;
		RECT	6.215 275.605 6.265 275.735 ;
		RECT	3.6 275.835 3.65 275.965 ;
		RECT	1.625 276.295 1.675 276.425 ;
		RECT	1.88 276.335 2.01 276.385 ;
		RECT	5.01 276.335 5.14 276.385 ;
		RECT	3.6 278.255 3.65 278.385 ;
		RECT	1.44 278.485 1.49 278.615 ;
		RECT	2.11 278.485 2.16 278.615 ;
		RECT	3.09 278.485 3.14 278.615 ;
		RECT	4.38 278.485 4.43 278.615 ;
		RECT	6.215 278.485 6.265 278.615 ;
		RECT	3.6 278.715 3.65 278.845 ;
		RECT	1.625 279.175 1.675 279.305 ;
		RECT	1.88 279.215 2.01 279.265 ;
		RECT	5.01 279.215 5.14 279.265 ;
		RECT	3.6 281.135 3.65 281.265 ;
		RECT	1.44 281.365 1.49 281.495 ;
		RECT	2.11 281.365 2.16 281.495 ;
		RECT	3.09 281.365 3.14 281.495 ;
		RECT	4.38 281.365 4.43 281.495 ;
		RECT	6.215 281.365 6.265 281.495 ;
		RECT	3.6 281.595 3.65 281.725 ;
		RECT	1.625 282.055 1.675 282.185 ;
		RECT	1.88 282.095 2.01 282.145 ;
		RECT	5.01 282.095 5.14 282.145 ;
		RECT	3.6 284.015 3.65 284.145 ;
		RECT	1.44 284.245 1.49 284.375 ;
		RECT	2.11 284.245 2.16 284.375 ;
		RECT	3.09 284.245 3.14 284.375 ;
		RECT	4.38 284.245 4.43 284.375 ;
		RECT	6.215 284.245 6.265 284.375 ;
		RECT	3.6 284.475 3.65 284.605 ;
		RECT	1.625 284.935 1.675 285.065 ;
		RECT	1.88 284.975 2.01 285.025 ;
		RECT	5.01 284.975 5.14 285.025 ;
		RECT	3.6 286.895 3.65 287.025 ;
		RECT	1.44 287.125 1.49 287.255 ;
		RECT	2.11 287.125 2.16 287.255 ;
		RECT	3.09 287.125 3.14 287.255 ;
		RECT	4.38 287.125 4.43 287.255 ;
		RECT	6.215 287.125 6.265 287.255 ;
		RECT	3.6 235.515 3.65 235.645 ;
		RECT	1.625 235.975 1.675 236.105 ;
		RECT	1.88 236.015 2.01 236.065 ;
		RECT	5.01 236.015 5.14 236.065 ;
		RECT	3.6 237.935 3.65 238.065 ;
		RECT	1.44 238.165 1.49 238.295 ;
		RECT	2.11 238.165 2.16 238.295 ;
		RECT	3.09 238.165 3.14 238.295 ;
		RECT	4.38 238.165 4.43 238.295 ;
		RECT	6.215 238.165 6.265 238.295 ;
		RECT	3.6 287.355 3.65 287.485 ;
		RECT	1.625 287.815 1.675 287.945 ;
		RECT	1.88 287.855 2.01 287.905 ;
		RECT	5.01 287.855 5.14 287.905 ;
		RECT	3.6 289.775 3.65 289.905 ;
		RECT	1.44 290.005 1.49 290.135 ;
		RECT	2.11 290.005 2.16 290.135 ;
		RECT	3.09 290.005 3.14 290.135 ;
		RECT	4.38 290.005 4.43 290.135 ;
		RECT	6.215 290.005 6.265 290.135 ;
		RECT	3.6 290.235 3.65 290.365 ;
		RECT	1.625 290.695 1.675 290.825 ;
		RECT	1.88 290.735 2.01 290.785 ;
		RECT	5.01 290.735 5.14 290.785 ;
		RECT	3.6 292.655 3.65 292.785 ;
		RECT	1.44 292.885 1.49 293.015 ;
		RECT	2.11 292.885 2.16 293.015 ;
		RECT	3.09 292.885 3.14 293.015 ;
		RECT	4.38 292.885 4.43 293.015 ;
		RECT	6.215 292.885 6.265 293.015 ;
		RECT	3.6 293.115 3.65 293.245 ;
		RECT	1.625 293.575 1.675 293.705 ;
		RECT	1.88 293.615 2.01 293.665 ;
		RECT	5.01 293.615 5.14 293.665 ;
		RECT	3.6 295.535 3.65 295.665 ;
		RECT	1.44 295.765 1.49 295.895 ;
		RECT	2.11 295.765 2.16 295.895 ;
		RECT	3.09 295.765 3.14 295.895 ;
		RECT	4.38 295.765 4.43 295.895 ;
		RECT	6.215 295.765 6.265 295.895 ;
		RECT	3.6 295.995 3.65 296.125 ;
		RECT	1.625 296.455 1.675 296.585 ;
		RECT	1.88 296.495 2.01 296.545 ;
		RECT	5.01 296.495 5.14 296.545 ;
		RECT	3.6 298.415 3.65 298.545 ;
		RECT	1.44 298.645 1.49 298.775 ;
		RECT	2.11 298.645 2.16 298.775 ;
		RECT	3.09 298.645 3.14 298.775 ;
		RECT	4.38 298.645 4.43 298.775 ;
		RECT	6.215 298.645 6.265 298.775 ;
		RECT	3.6 298.875 3.65 299.005 ;
		RECT	1.625 299.335 1.675 299.465 ;
		RECT	1.88 299.375 2.01 299.425 ;
		RECT	5.01 299.375 5.14 299.425 ;
		RECT	3.6 301.295 3.65 301.425 ;
		RECT	1.44 301.525 1.49 301.655 ;
		RECT	2.11 301.525 2.16 301.655 ;
		RECT	3.09 301.525 3.14 301.655 ;
		RECT	4.38 301.525 4.43 301.655 ;
		RECT	6.215 301.525 6.265 301.655 ;
		RECT	3.6 301.755 3.65 301.885 ;
		RECT	1.625 302.215 1.675 302.345 ;
		RECT	1.88 302.255 2.01 302.305 ;
		RECT	5.01 302.255 5.14 302.305 ;
		RECT	3.6 304.175 3.65 304.305 ;
		RECT	1.44 304.405 1.49 304.535 ;
		RECT	2.11 304.405 2.16 304.535 ;
		RECT	3.09 304.405 3.14 304.535 ;
		RECT	4.38 304.405 4.43 304.535 ;
		RECT	6.215 304.405 6.265 304.535 ;
		RECT	3.6 304.635 3.65 304.765 ;
		RECT	1.625 305.095 1.675 305.225 ;
		RECT	1.88 305.135 2.01 305.185 ;
		RECT	5.01 305.135 5.14 305.185 ;
		RECT	3.6 307.055 3.65 307.185 ;
		RECT	1.44 307.285 1.49 307.415 ;
		RECT	2.11 307.285 2.16 307.415 ;
		RECT	3.09 307.285 3.14 307.415 ;
		RECT	4.38 307.285 4.43 307.415 ;
		RECT	6.215 307.285 6.265 307.415 ;
		RECT	3.6 307.515 3.65 307.645 ;
		RECT	1.625 307.975 1.675 308.105 ;
		RECT	1.88 308.015 2.01 308.065 ;
		RECT	5.01 308.015 5.14 308.065 ;
		RECT	3.6 309.935 3.65 310.065 ;
		RECT	1.44 310.165 1.49 310.295 ;
		RECT	2.11 310.165 2.16 310.295 ;
		RECT	3.09 310.165 3.14 310.295 ;
		RECT	4.38 310.165 4.43 310.295 ;
		RECT	6.215 310.165 6.265 310.295 ;
		RECT	3.6 310.395 3.65 310.525 ;
		RECT	1.625 310.855 1.675 310.985 ;
		RECT	1.88 310.895 2.01 310.945 ;
		RECT	5.01 310.895 5.14 310.945 ;
		RECT	3.6 312.815 3.65 312.945 ;
		RECT	1.44 313.045 1.49 313.175 ;
		RECT	2.11 313.045 2.16 313.175 ;
		RECT	3.09 313.045 3.14 313.175 ;
		RECT	4.38 313.045 4.43 313.175 ;
		RECT	6.215 313.045 6.265 313.175 ;
		RECT	3.6 313.275 3.65 313.405 ;
		RECT	1.625 313.735 1.675 313.865 ;
		RECT	1.88 313.775 2.01 313.825 ;
		RECT	5.01 313.775 5.14 313.825 ;
		RECT	3.6 315.695 3.65 315.825 ;
		RECT	1.44 315.925 1.49 316.055 ;
		RECT	2.11 315.925 2.16 316.055 ;
		RECT	3.09 315.925 3.14 316.055 ;
		RECT	4.38 315.925 4.43 316.055 ;
		RECT	6.215 315.925 6.265 316.055 ;
		RECT	3.6 238.395 3.65 238.525 ;
		RECT	1.625 238.855 1.675 238.985 ;
		RECT	1.88 238.895 2.01 238.945 ;
		RECT	5.01 238.895 5.14 238.945 ;
		RECT	3.6 240.815 3.65 240.945 ;
		RECT	1.44 241.045 1.49 241.175 ;
		RECT	2.11 241.045 2.16 241.175 ;
		RECT	3.09 241.045 3.14 241.175 ;
		RECT	4.38 241.045 4.43 241.175 ;
		RECT	6.215 241.045 6.265 241.175 ;
		RECT	3.6 316.155 3.65 316.285 ;
		RECT	1.625 316.615 1.675 316.745 ;
		RECT	1.88 316.655 2.01 316.705 ;
		RECT	5.01 316.655 5.14 316.705 ;
		RECT	3.6 318.575 3.65 318.705 ;
		RECT	1.44 318.805 1.49 318.935 ;
		RECT	2.11 318.805 2.16 318.935 ;
		RECT	3.09 318.805 3.14 318.935 ;
		RECT	4.38 318.805 4.43 318.935 ;
		RECT	6.215 318.805 6.265 318.935 ;
		RECT	3.6 319.035 3.65 319.165 ;
		RECT	1.625 319.495 1.675 319.625 ;
		RECT	1.88 319.535 2.01 319.585 ;
		RECT	5.01 319.535 5.14 319.585 ;
		RECT	3.6 321.455 3.65 321.585 ;
		RECT	1.44 321.685 1.49 321.815 ;
		RECT	2.11 321.685 2.16 321.815 ;
		RECT	3.09 321.685 3.14 321.815 ;
		RECT	4.38 321.685 4.43 321.815 ;
		RECT	6.215 321.685 6.265 321.815 ;
		RECT	3.6 321.915 3.65 322.045 ;
		RECT	1.625 322.375 1.675 322.505 ;
		RECT	1.88 322.415 2.01 322.465 ;
		RECT	5.01 322.415 5.14 322.465 ;
		RECT	3.6 324.335 3.65 324.465 ;
		RECT	1.44 324.565 1.49 324.695 ;
		RECT	2.11 324.565 2.16 324.695 ;
		RECT	3.09 324.565 3.14 324.695 ;
		RECT	4.38 324.565 4.43 324.695 ;
		RECT	6.215 324.565 6.265 324.695 ;
		RECT	3.6 324.795 3.65 324.925 ;
		RECT	1.625 325.255 1.675 325.385 ;
		RECT	1.88 325.295 2.01 325.345 ;
		RECT	5.01 325.295 5.14 325.345 ;
		RECT	3.6 327.215 3.65 327.345 ;
		RECT	1.44 327.445 1.49 327.575 ;
		RECT	2.11 327.445 2.16 327.575 ;
		RECT	3.09 327.445 3.14 327.575 ;
		RECT	4.38 327.445 4.43 327.575 ;
		RECT	6.215 327.445 6.265 327.575 ;
		RECT	3.6 327.675 3.65 327.805 ;
		RECT	1.625 328.135 1.675 328.265 ;
		RECT	1.88 328.175 2.01 328.225 ;
		RECT	5.01 328.175 5.14 328.225 ;
		RECT	3.6 330.095 3.65 330.225 ;
		RECT	1.44 330.325 1.49 330.455 ;
		RECT	2.11 330.325 2.16 330.455 ;
		RECT	3.09 330.325 3.14 330.455 ;
		RECT	4.38 330.325 4.43 330.455 ;
		RECT	6.215 330.325 6.265 330.455 ;
		RECT	3.6 330.555 3.65 330.685 ;
		RECT	1.625 331.015 1.675 331.145 ;
		RECT	1.88 331.055 2.01 331.105 ;
		RECT	5.01 331.055 5.14 331.105 ;
		RECT	3.6 332.975 3.65 333.105 ;
		RECT	1.44 333.205 1.49 333.335 ;
		RECT	2.11 333.205 2.16 333.335 ;
		RECT	3.09 333.205 3.14 333.335 ;
		RECT	4.38 333.205 4.43 333.335 ;
		RECT	6.215 333.205 6.265 333.335 ;
		RECT	3.6 333.435 3.65 333.565 ;
		RECT	1.625 333.895 1.675 334.025 ;
		RECT	1.88 333.935 2.01 333.985 ;
		RECT	5.01 333.935 5.14 333.985 ;
		RECT	3.6 335.855 3.65 335.985 ;
		RECT	1.44 336.085 1.49 336.215 ;
		RECT	2.11 336.085 2.16 336.215 ;
		RECT	3.09 336.085 3.14 336.215 ;
		RECT	4.38 336.085 4.43 336.215 ;
		RECT	6.215 336.085 6.265 336.215 ;
		RECT	3.6 336.315 3.65 336.445 ;
		RECT	1.625 336.775 1.675 336.905 ;
		RECT	1.88 336.815 2.01 336.865 ;
		RECT	5.01 336.815 5.14 336.865 ;
		RECT	3.6 338.735 3.65 338.865 ;
		RECT	1.44 338.965 1.49 339.095 ;
		RECT	2.11 338.965 2.16 339.095 ;
		RECT	3.09 338.965 3.14 339.095 ;
		RECT	4.38 338.965 4.43 339.095 ;
		RECT	6.215 338.965 6.265 339.095 ;
		RECT	3.6 339.195 3.65 339.325 ;
		RECT	1.625 339.655 1.675 339.785 ;
		RECT	1.88 339.695 2.01 339.745 ;
		RECT	5.01 339.695 5.14 339.745 ;
		RECT	3.6 341.615 3.65 341.745 ;
		RECT	1.44 341.845 1.49 341.975 ;
		RECT	2.11 341.845 2.16 341.975 ;
		RECT	3.09 341.845 3.14 341.975 ;
		RECT	4.38 341.845 4.43 341.975 ;
		RECT	6.215 341.845 6.265 341.975 ;
		RECT	3.6 342.075 3.65 342.205 ;
		RECT	1.625 342.535 1.675 342.665 ;
		RECT	1.88 342.575 2.01 342.625 ;
		RECT	5.01 342.575 5.14 342.625 ;
		RECT	3.6 344.495 3.65 344.625 ;
		RECT	1.44 344.725 1.49 344.855 ;
		RECT	2.11 344.725 2.16 344.855 ;
		RECT	3.09 344.725 3.14 344.855 ;
		RECT	4.38 344.725 4.43 344.855 ;
		RECT	6.215 344.725 6.265 344.855 ;
		RECT	3.6 241.275 3.65 241.405 ;
		RECT	1.625 241.735 1.675 241.865 ;
		RECT	1.88 241.775 2.01 241.825 ;
		RECT	5.01 241.775 5.14 241.825 ;
		RECT	3.6 243.695 3.65 243.825 ;
		RECT	1.44 243.925 1.49 244.055 ;
		RECT	2.11 243.925 2.16 244.055 ;
		RECT	3.09 243.925 3.14 244.055 ;
		RECT	4.38 243.925 4.43 244.055 ;
		RECT	6.215 243.925 6.265 244.055 ;
		RECT	3.6 344.955 3.65 345.085 ;
		RECT	1.625 345.415 1.675 345.545 ;
		RECT	1.88 345.455 2.01 345.505 ;
		RECT	5.01 345.455 5.14 345.505 ;
		RECT	3.6 347.375 3.65 347.505 ;
		RECT	1.44 347.605 1.49 347.735 ;
		RECT	2.11 347.605 2.16 347.735 ;
		RECT	3.09 347.605 3.14 347.735 ;
		RECT	4.38 347.605 4.43 347.735 ;
		RECT	6.215 347.605 6.265 347.735 ;
		RECT	3.6 347.835 3.65 347.965 ;
		RECT	1.625 348.295 1.675 348.425 ;
		RECT	1.88 348.335 2.01 348.385 ;
		RECT	5.01 348.335 5.14 348.385 ;
		RECT	3.6 350.255 3.65 350.385 ;
		RECT	1.44 350.485 1.49 350.615 ;
		RECT	2.11 350.485 2.16 350.615 ;
		RECT	3.09 350.485 3.14 350.615 ;
		RECT	4.38 350.485 4.43 350.615 ;
		RECT	6.215 350.485 6.265 350.615 ;
		RECT	3.6 350.715 3.65 350.845 ;
		RECT	1.625 351.175 1.675 351.305 ;
		RECT	1.88 351.215 2.01 351.265 ;
		RECT	5.01 351.215 5.14 351.265 ;
		RECT	3.6 353.135 3.65 353.265 ;
		RECT	1.44 353.365 1.49 353.495 ;
		RECT	2.11 353.365 2.16 353.495 ;
		RECT	3.09 353.365 3.14 353.495 ;
		RECT	4.38 353.365 4.43 353.495 ;
		RECT	6.215 353.365 6.265 353.495 ;
		RECT	3.6 353.595 3.65 353.725 ;
		RECT	1.625 354.055 1.675 354.185 ;
		RECT	1.88 354.095 2.01 354.145 ;
		RECT	5.01 354.095 5.14 354.145 ;
		RECT	3.6 356.015 3.65 356.145 ;
		RECT	1.44 356.245 1.49 356.375 ;
		RECT	2.11 356.245 2.16 356.375 ;
		RECT	3.09 356.245 3.14 356.375 ;
		RECT	4.38 356.245 4.43 356.375 ;
		RECT	6.215 356.245 6.265 356.375 ;
		RECT	3.6 356.475 3.65 356.605 ;
		RECT	1.625 356.935 1.675 357.065 ;
		RECT	1.88 356.975 2.01 357.025 ;
		RECT	5.01 356.975 5.14 357.025 ;
		RECT	3.6 358.895 3.65 359.025 ;
		RECT	1.44 359.125 1.49 359.255 ;
		RECT	2.11 359.125 2.16 359.255 ;
		RECT	3.09 359.125 3.14 359.255 ;
		RECT	4.38 359.125 4.43 359.255 ;
		RECT	6.215 359.125 6.265 359.255 ;
		RECT	3.6 359.355 3.65 359.485 ;
		RECT	1.625 359.815 1.675 359.945 ;
		RECT	1.88 359.855 2.01 359.905 ;
		RECT	5.01 359.855 5.14 359.905 ;
		RECT	3.6 361.775 3.65 361.905 ;
		RECT	1.44 362.005 1.49 362.135 ;
		RECT	2.11 362.005 2.16 362.135 ;
		RECT	3.09 362.005 3.14 362.135 ;
		RECT	4.38 362.005 4.43 362.135 ;
		RECT	6.215 362.005 6.265 362.135 ;
		RECT	3.6 362.235 3.65 362.365 ;
		RECT	1.625 362.695 1.675 362.825 ;
		RECT	1.88 362.735 2.01 362.785 ;
		RECT	5.01 362.735 5.14 362.785 ;
		RECT	3.6 364.655 3.65 364.785 ;
		RECT	1.44 364.885 1.49 365.015 ;
		RECT	2.11 364.885 2.16 365.015 ;
		RECT	3.09 364.885 3.14 365.015 ;
		RECT	4.38 364.885 4.43 365.015 ;
		RECT	6.215 364.885 6.265 365.015 ;
		RECT	3.6 365.115 3.65 365.245 ;
		RECT	1.625 365.575 1.675 365.705 ;
		RECT	1.88 365.615 2.01 365.665 ;
		RECT	5.01 365.615 5.14 365.665 ;
		RECT	3.6 367.535 3.65 367.665 ;
		RECT	1.44 367.765 1.49 367.895 ;
		RECT	2.11 367.765 2.16 367.895 ;
		RECT	3.09 367.765 3.14 367.895 ;
		RECT	4.38 367.765 4.43 367.895 ;
		RECT	6.215 367.765 6.265 367.895 ;
		RECT	3.6 367.995 3.65 368.125 ;
		RECT	1.625 368.455 1.675 368.585 ;
		RECT	1.88 368.495 2.01 368.545 ;
		RECT	5.01 368.495 5.14 368.545 ;
		RECT	3.6 370.415 3.65 370.545 ;
		RECT	1.44 370.645 1.49 370.775 ;
		RECT	2.11 370.645 2.16 370.775 ;
		RECT	3.09 370.645 3.14 370.775 ;
		RECT	4.38 370.645 4.43 370.775 ;
		RECT	6.215 370.645 6.265 370.775 ;
		RECT	3.6 370.875 3.65 371.005 ;
		RECT	1.625 371.335 1.675 371.465 ;
		RECT	1.88 371.375 2.01 371.425 ;
		RECT	5.01 371.375 5.14 371.425 ;
		RECT	3.6 373.295 3.65 373.425 ;
		RECT	1.44 373.525 1.49 373.655 ;
		RECT	2.11 373.525 2.16 373.655 ;
		RECT	3.09 373.525 3.14 373.655 ;
		RECT	4.38 373.525 4.43 373.655 ;
		RECT	6.215 373.525 6.265 373.655 ;
		RECT	3.6 244.155 3.65 244.285 ;
		RECT	1.625 244.615 1.675 244.745 ;
		RECT	1.88 244.655 2.01 244.705 ;
		RECT	5.01 244.655 5.14 244.705 ;
		RECT	3.6 246.575 3.65 246.705 ;
		RECT	1.44 246.805 1.49 246.935 ;
		RECT	2.11 246.805 2.16 246.935 ;
		RECT	3.09 246.805 3.14 246.935 ;
		RECT	4.38 246.805 4.43 246.935 ;
		RECT	6.215 246.805 6.265 246.935 ;
		RECT	3.6 373.755 3.65 373.885 ;
		RECT	1.625 374.215 1.675 374.345 ;
		RECT	1.88 374.255 2.01 374.305 ;
		RECT	5.01 374.255 5.14 374.305 ;
		RECT	3.6 376.175 3.65 376.305 ;
		RECT	1.44 376.405 1.49 376.535 ;
		RECT	2.11 376.405 2.16 376.535 ;
		RECT	3.09 376.405 3.14 376.535 ;
		RECT	4.38 376.405 4.43 376.535 ;
		RECT	6.215 376.405 6.265 376.535 ;
		RECT	3.6 376.635 3.65 376.765 ;
		RECT	1.625 377.095 1.675 377.225 ;
		RECT	1.88 377.135 2.01 377.185 ;
		RECT	5.01 377.135 5.14 377.185 ;
		RECT	3.6 379.055 3.65 379.185 ;
		RECT	1.44 379.285 1.49 379.415 ;
		RECT	2.11 379.285 2.16 379.415 ;
		RECT	3.09 379.285 3.14 379.415 ;
		RECT	4.38 379.285 4.43 379.415 ;
		RECT	6.215 379.285 6.265 379.415 ;
		RECT	3.6 379.515 3.65 379.645 ;
		RECT	1.625 379.975 1.675 380.105 ;
		RECT	1.88 380.015 2.01 380.065 ;
		RECT	5.01 380.015 5.14 380.065 ;
		RECT	3.6 381.935 3.65 382.065 ;
		RECT	1.44 382.165 1.49 382.295 ;
		RECT	2.11 382.165 2.16 382.295 ;
		RECT	3.09 382.165 3.14 382.295 ;
		RECT	4.38 382.165 4.43 382.295 ;
		RECT	6.215 382.165 6.265 382.295 ;
		RECT	3.6 382.395 3.65 382.525 ;
		RECT	1.625 382.855 1.675 382.985 ;
		RECT	1.88 382.895 2.01 382.945 ;
		RECT	5.01 382.895 5.14 382.945 ;
		RECT	3.6 384.815 3.65 384.945 ;
		RECT	1.44 385.045 1.49 385.175 ;
		RECT	2.11 385.045 2.16 385.175 ;
		RECT	3.09 385.045 3.14 385.175 ;
		RECT	4.38 385.045 4.43 385.175 ;
		RECT	6.215 385.045 6.265 385.175 ;
		RECT	3.6 385.275 3.65 385.405 ;
		RECT	1.625 385.735 1.675 385.865 ;
		RECT	1.88 385.775 2.01 385.825 ;
		RECT	5.01 385.775 5.14 385.825 ;
		RECT	3.6 387.695 3.65 387.825 ;
		RECT	1.44 387.925 1.49 388.055 ;
		RECT	2.11 387.925 2.16 388.055 ;
		RECT	3.09 387.925 3.14 388.055 ;
		RECT	4.38 387.925 4.43 388.055 ;
		RECT	6.215 387.925 6.265 388.055 ;
		RECT	3.6 388.155 3.65 388.285 ;
		RECT	1.625 388.615 1.675 388.745 ;
		RECT	1.88 388.655 2.01 388.705 ;
		RECT	5.01 388.655 5.14 388.705 ;
		RECT	3.6 390.575 3.65 390.705 ;
		RECT	1.44 390.805 1.49 390.935 ;
		RECT	2.11 390.805 2.16 390.935 ;
		RECT	3.09 390.805 3.14 390.935 ;
		RECT	4.38 390.805 4.43 390.935 ;
		RECT	6.215 390.805 6.265 390.935 ;
		RECT	3.6 391.035 3.65 391.165 ;
		RECT	1.625 391.495 1.675 391.625 ;
		RECT	1.88 391.535 2.01 391.585 ;
		RECT	5.01 391.535 5.14 391.585 ;
		RECT	3.6 393.455 3.65 393.585 ;
		RECT	1.44 393.685 1.49 393.815 ;
		RECT	2.11 393.685 2.16 393.815 ;
		RECT	3.09 393.685 3.14 393.815 ;
		RECT	4.38 393.685 4.43 393.815 ;
		RECT	6.215 393.685 6.265 393.815 ;
		RECT	3.6 393.915 3.65 394.045 ;
		RECT	1.625 394.375 1.675 394.505 ;
		RECT	1.88 394.415 2.01 394.465 ;
		RECT	5.01 394.415 5.14 394.465 ;
		RECT	3.6 396.335 3.65 396.465 ;
		RECT	1.44 396.565 1.49 396.695 ;
		RECT	2.11 396.565 2.16 396.695 ;
		RECT	3.09 396.565 3.14 396.695 ;
		RECT	4.38 396.565 4.43 396.695 ;
		RECT	6.215 396.565 6.265 396.695 ;
		RECT	3.6 396.795 3.65 396.925 ;
		RECT	1.625 397.255 1.675 397.385 ;
		RECT	1.88 397.295 2.01 397.345 ;
		RECT	5.01 397.295 5.14 397.345 ;
		RECT	3.6 399.215 3.65 399.345 ;
		RECT	1.44 399.445 1.49 399.575 ;
		RECT	2.11 399.445 2.16 399.575 ;
		RECT	3.09 399.445 3.14 399.575 ;
		RECT	4.38 399.445 4.43 399.575 ;
		RECT	6.215 399.445 6.265 399.575 ;
		RECT	3.6 399.675 3.65 399.805 ;
		RECT	1.625 400.135 1.675 400.265 ;
		RECT	1.88 400.175 2.01 400.225 ;
		RECT	5.01 400.175 5.14 400.225 ;
		RECT	3.6 402.095 3.65 402.225 ;
		RECT	1.44 402.325 1.49 402.455 ;
		RECT	2.11 402.325 2.16 402.455 ;
		RECT	3.09 402.325 3.14 402.455 ;
		RECT	4.38 402.325 4.43 402.455 ;
		RECT	6.215 402.325 6.265 402.455 ;
		RECT	3.6 247.035 3.65 247.165 ;
		RECT	1.625 247.495 1.675 247.625 ;
		RECT	1.88 247.535 2.01 247.585 ;
		RECT	5.01 247.535 5.14 247.585 ;
		RECT	3.6 249.455 3.65 249.585 ;
		RECT	1.44 249.685 1.49 249.815 ;
		RECT	2.11 249.685 2.16 249.815 ;
		RECT	3.09 249.685 3.14 249.815 ;
		RECT	4.38 249.685 4.43 249.815 ;
		RECT	6.215 249.685 6.265 249.815 ;
		RECT	3.6 402.555 3.65 402.685 ;
		RECT	1.625 403.015 1.675 403.145 ;
		RECT	1.88 403.055 2.01 403.105 ;
		RECT	5.01 403.055 5.14 403.105 ;
		RECT	3.6 404.975 3.65 405.105 ;
		RECT	1.44 405.205 1.49 405.335 ;
		RECT	2.11 405.205 2.16 405.335 ;
		RECT	3.09 405.205 3.14 405.335 ;
		RECT	4.38 405.205 4.43 405.335 ;
		RECT	6.215 405.205 6.265 405.335 ;
		RECT	3.6 405.435 3.65 405.565 ;
		RECT	1.625 405.895 1.675 406.025 ;
		RECT	1.88 405.935 2.01 405.985 ;
		RECT	5.01 405.935 5.14 405.985 ;
		RECT	3.6 407.855 3.65 407.985 ;
		RECT	1.44 408.085 1.49 408.215 ;
		RECT	2.11 408.085 2.16 408.215 ;
		RECT	3.09 408.085 3.14 408.215 ;
		RECT	4.38 408.085 4.43 408.215 ;
		RECT	6.215 408.085 6.265 408.215 ;
		RECT	3.6 408.315 3.65 408.445 ;
		RECT	1.625 408.775 1.675 408.905 ;
		RECT	1.88 408.815 2.01 408.865 ;
		RECT	5.01 408.815 5.14 408.865 ;
		RECT	3.6 410.735 3.65 410.865 ;
		RECT	1.44 410.965 1.49 411.095 ;
		RECT	2.11 410.965 2.16 411.095 ;
		RECT	3.09 410.965 3.14 411.095 ;
		RECT	4.38 410.965 4.43 411.095 ;
		RECT	6.215 410.965 6.265 411.095 ;
		RECT	3.6 249.915 3.65 250.045 ;
		RECT	1.625 250.375 1.675 250.505 ;
		RECT	1.88 250.415 2.01 250.465 ;
		RECT	5.01 250.415 5.14 250.465 ;
		RECT	3.6 252.335 3.65 252.465 ;
		RECT	1.44 252.565 1.49 252.695 ;
		RECT	2.11 252.565 2.16 252.695 ;
		RECT	3.09 252.565 3.14 252.695 ;
		RECT	4.38 252.565 4.43 252.695 ;
		RECT	6.215 252.565 6.265 252.695 ;
		RECT	3.6 252.795 3.65 252.925 ;
		RECT	1.625 253.255 1.675 253.385 ;
		RECT	1.88 253.295 2.01 253.345 ;
		RECT	5.01 253.295 5.14 253.345 ;
		RECT	3.6 255.215 3.65 255.345 ;
		RECT	1.44 255.445 1.49 255.575 ;
		RECT	2.11 255.445 2.16 255.575 ;
		RECT	3.09 255.445 3.14 255.575 ;
		RECT	4.38 255.445 4.43 255.575 ;
		RECT	6.215 255.445 6.265 255.575 ;
		RECT	3.6 255.675 3.65 255.805 ;
		RECT	1.625 256.135 1.675 256.265 ;
		RECT	1.88 256.175 2.01 256.225 ;
		RECT	5.01 256.175 5.14 256.225 ;
		RECT	3.6 258.095 3.65 258.225 ;
		RECT	1.44 258.325 1.49 258.455 ;
		RECT	2.11 258.325 2.16 258.455 ;
		RECT	3.09 258.325 3.14 258.455 ;
		RECT	4.38 258.325 4.43 258.455 ;
		RECT	6.215 258.325 6.265 258.455 ;
		RECT	3.6 411.195 3.65 411.325 ;
		RECT	1.625 411.655 1.675 411.785 ;
		RECT	1.88 411.695 2.01 411.745 ;
		RECT	5.01 411.695 5.14 411.745 ;
		RECT	3.6 413.615 3.65 413.745 ;
		RECT	1.44 413.845 1.49 413.975 ;
		RECT	2.11 413.845 2.16 413.975 ;
		RECT	3.09 413.845 3.14 413.975 ;
		RECT	4.38 413.845 4.43 413.975 ;
		RECT	6.215 413.845 6.265 413.975 ;
		RECT	3.6 229.755 3.65 229.885 ;
		RECT	1.625 230.215 1.675 230.345 ;
		RECT	1.88 230.255 2.01 230.305 ;
		RECT	5.01 230.255 5.14 230.305 ;
		RECT	3.6 232.175 3.65 232.305 ;
		RECT	1.44 232.405 1.49 232.535 ;
		RECT	2.11 232.405 2.16 232.535 ;
		RECT	3.09 232.405 3.14 232.535 ;
		RECT	4.38 232.405 4.43 232.535 ;
		RECT	6.215 232.405 6.265 232.535 ;
		RECT	0.435 230.215 0.485 230.345 ;
		RECT	0.435 229.755 0.485 229.885 ;
		RECT	0.435 232.175 0.485 232.305 ;
		RECT	0.435 233.095 0.485 233.225 ;
		RECT	0.435 232.635 0.485 232.765 ;
		RECT	0.435 235.055 0.485 235.185 ;
		RECT	0.435 259.015 0.485 259.145 ;
		RECT	0.435 258.555 0.485 258.685 ;
		RECT	0.435 260.975 0.485 261.105 ;
		RECT	0.435 261.895 0.485 262.025 ;
		RECT	0.435 261.435 0.485 261.565 ;
		RECT	0.435 263.855 0.485 263.985 ;
		RECT	0.435 264.775 0.485 264.905 ;
		RECT	0.435 264.315 0.485 264.445 ;
		RECT	0.435 266.735 0.485 266.865 ;
		RECT	0.435 267.655 0.485 267.785 ;
		RECT	0.435 267.195 0.485 267.325 ;
		RECT	0.435 269.615 0.485 269.745 ;
		RECT	0.435 270.535 0.485 270.665 ;
		RECT	0.435 270.075 0.485 270.205 ;
		RECT	0.435 272.495 0.485 272.625 ;
		RECT	0.435 273.415 0.485 273.545 ;
		RECT	0.435 272.955 0.485 273.085 ;
		RECT	0.435 275.375 0.485 275.505 ;
		RECT	0.435 276.295 0.485 276.425 ;
		RECT	0.435 275.835 0.485 275.965 ;
		RECT	0.435 278.255 0.485 278.385 ;
		RECT	0.435 279.175 0.485 279.305 ;
		RECT	0.435 278.715 0.485 278.845 ;
		RECT	0.435 281.135 0.485 281.265 ;
		RECT	0.435 282.055 0.485 282.185 ;
		RECT	0.435 281.595 0.485 281.725 ;
		RECT	0.435 284.015 0.485 284.145 ;
		RECT	0.435 284.935 0.485 285.065 ;
		RECT	0.435 284.475 0.485 284.605 ;
		RECT	0.435 286.895 0.485 287.025 ;
		RECT	0.435 235.975 0.485 236.105 ;
		RECT	0.435 235.515 0.485 235.645 ;
		RECT	0.435 237.935 0.485 238.065 ;
		RECT	0.435 287.815 0.485 287.945 ;
		RECT	0.435 287.355 0.485 287.485 ;
		RECT	0.435 289.775 0.485 289.905 ;
		RECT	0.435 290.695 0.485 290.825 ;
		RECT	0.435 290.235 0.485 290.365 ;
		RECT	0.435 292.655 0.485 292.785 ;
		RECT	0.435 293.575 0.485 293.705 ;
		RECT	0.435 293.115 0.485 293.245 ;
		RECT	0.435 295.535 0.485 295.665 ;
		RECT	0.435 296.455 0.485 296.585 ;
		RECT	0.435 295.995 0.485 296.125 ;
		RECT	0.435 298.415 0.485 298.545 ;
		RECT	0.435 299.335 0.485 299.465 ;
		RECT	0.435 298.875 0.485 299.005 ;
		RECT	0.435 301.295 0.485 301.425 ;
		RECT	0.435 302.215 0.485 302.345 ;
		RECT	0.435 301.755 0.485 301.885 ;
		RECT	0.435 304.175 0.485 304.305 ;
		RECT	0.435 305.095 0.485 305.225 ;
		RECT	0.435 304.635 0.485 304.765 ;
		RECT	0.435 307.055 0.485 307.185 ;
		RECT	0.435 307.975 0.485 308.105 ;
		RECT	0.435 307.515 0.485 307.645 ;
		RECT	0.435 309.935 0.485 310.065 ;
		RECT	0.435 310.855 0.485 310.985 ;
		RECT	0.435 310.395 0.485 310.525 ;
		RECT	0.435 312.815 0.485 312.945 ;
		RECT	0.435 313.735 0.485 313.865 ;
		RECT	0.435 313.275 0.485 313.405 ;
		RECT	0.435 315.695 0.485 315.825 ;
		RECT	0.435 238.855 0.485 238.985 ;
		RECT	0.435 238.395 0.485 238.525 ;
		RECT	0.435 240.815 0.485 240.945 ;
		RECT	0.435 316.615 0.485 316.745 ;
		RECT	0.435 316.155 0.485 316.285 ;
		RECT	0.435 318.575 0.485 318.705 ;
		RECT	0.435 319.495 0.485 319.625 ;
		RECT	0.435 319.035 0.485 319.165 ;
		RECT	0.435 321.455 0.485 321.585 ;
		RECT	0.435 322.375 0.485 322.505 ;
		RECT	0.435 321.915 0.485 322.045 ;
		RECT	0.435 324.335 0.485 324.465 ;
		RECT	0.435 325.255 0.485 325.385 ;
		RECT	0.435 324.795 0.485 324.925 ;
		RECT	0.435 327.215 0.485 327.345 ;
		RECT	0.435 328.135 0.485 328.265 ;
		RECT	0.435 327.675 0.485 327.805 ;
		RECT	0.435 330.095 0.485 330.225 ;
		RECT	0.435 331.015 0.485 331.145 ;
		RECT	0.435 330.555 0.485 330.685 ;
		RECT	0.435 332.975 0.485 333.105 ;
		RECT	0.435 333.895 0.485 334.025 ;
		RECT	0.435 333.435 0.485 333.565 ;
		RECT	0.435 335.855 0.485 335.985 ;
		RECT	0.435 336.775 0.485 336.905 ;
		RECT	0.435 336.315 0.485 336.445 ;
		RECT	0.435 338.735 0.485 338.865 ;
		RECT	0.435 339.655 0.485 339.785 ;
		RECT	0.435 339.195 0.485 339.325 ;
		RECT	0.435 341.615 0.485 341.745 ;
		RECT	0.435 342.535 0.485 342.665 ;
		RECT	0.435 342.075 0.485 342.205 ;
		RECT	0.435 344.495 0.485 344.625 ;
		RECT	0.435 241.735 0.485 241.865 ;
		RECT	0.435 241.275 0.485 241.405 ;
		RECT	0.435 243.695 0.485 243.825 ;
		RECT	0.435 345.415 0.485 345.545 ;
		RECT	0.435 344.955 0.485 345.085 ;
		RECT	0.435 347.375 0.485 347.505 ;
		RECT	0.435 348.295 0.485 348.425 ;
		RECT	0.435 347.835 0.485 347.965 ;
		RECT	0.435 350.255 0.485 350.385 ;
		RECT	0.435 351.175 0.485 351.305 ;
		RECT	0.435 350.715 0.485 350.845 ;
		RECT	0.435 353.135 0.485 353.265 ;
		RECT	0.435 354.055 0.485 354.185 ;
		RECT	0.435 353.595 0.485 353.725 ;
		RECT	0.435 356.015 0.485 356.145 ;
		RECT	0.435 356.935 0.485 357.065 ;
		RECT	0.435 356.475 0.485 356.605 ;
		RECT	0.435 358.895 0.485 359.025 ;
		RECT	0.435 359.815 0.485 359.945 ;
		RECT	0.435 359.355 0.485 359.485 ;
		RECT	0.435 361.775 0.485 361.905 ;
		RECT	0.435 362.695 0.485 362.825 ;
		RECT	0.435 362.235 0.485 362.365 ;
		RECT	0.435 364.655 0.485 364.785 ;
		RECT	0.435 365.575 0.485 365.705 ;
		RECT	0.435 365.115 0.485 365.245 ;
		RECT	0.435 367.535 0.485 367.665 ;
		RECT	0.435 368.455 0.485 368.585 ;
		RECT	0.435 367.995 0.485 368.125 ;
		RECT	0.435 370.415 0.485 370.545 ;
		RECT	0.435 371.335 0.485 371.465 ;
		RECT	0.435 370.875 0.485 371.005 ;
		RECT	0.435 373.295 0.485 373.425 ;
		RECT	0.435 244.615 0.485 244.745 ;
		RECT	0.435 244.155 0.485 244.285 ;
		RECT	0.435 246.575 0.485 246.705 ;
		RECT	0.435 374.215 0.485 374.345 ;
		RECT	0.435 373.755 0.485 373.885 ;
		RECT	0.435 376.175 0.485 376.305 ;
		RECT	0.435 377.095 0.485 377.225 ;
		RECT	0.435 376.635 0.485 376.765 ;
		RECT	0.435 379.055 0.485 379.185 ;
		RECT	0.435 379.975 0.485 380.105 ;
		RECT	0.435 379.515 0.485 379.645 ;
		RECT	0.435 381.935 0.485 382.065 ;
		RECT	0.435 382.855 0.485 382.985 ;
		RECT	0.435 382.395 0.485 382.525 ;
		RECT	0.435 384.815 0.485 384.945 ;
		RECT	0.435 385.735 0.485 385.865 ;
		RECT	0.435 385.275 0.485 385.405 ;
		RECT	0.435 387.695 0.485 387.825 ;
		RECT	0.435 388.615 0.485 388.745 ;
		RECT	0.435 388.155 0.485 388.285 ;
		RECT	0.435 390.575 0.485 390.705 ;
		RECT	0.435 391.495 0.485 391.625 ;
		RECT	0.435 391.035 0.485 391.165 ;
		RECT	0.435 393.455 0.485 393.585 ;
		RECT	0.435 394.375 0.485 394.505 ;
		RECT	0.435 393.915 0.485 394.045 ;
		RECT	0.435 396.335 0.485 396.465 ;
		RECT	0.435 397.255 0.485 397.385 ;
		RECT	0.435 396.795 0.485 396.925 ;
		RECT	0.435 399.215 0.485 399.345 ;
		RECT	0.435 400.135 0.485 400.265 ;
		RECT	0.435 399.675 0.485 399.805 ;
		RECT	0.435 402.095 0.485 402.225 ;
		RECT	0.435 247.495 0.485 247.625 ;
		RECT	0.435 247.035 0.485 247.165 ;
		RECT	0.435 249.455 0.485 249.585 ;
		RECT	0.435 403.015 0.485 403.145 ;
		RECT	0.435 402.555 0.485 402.685 ;
		RECT	0.435 404.975 0.485 405.105 ;
		RECT	0.435 405.895 0.485 406.025 ;
		RECT	0.435 405.435 0.485 405.565 ;
		RECT	0.435 407.855 0.485 407.985 ;
		RECT	0.435 408.775 0.485 408.905 ;
		RECT	0.435 408.315 0.485 408.445 ;
		RECT	0.435 410.735 0.485 410.865 ;
		RECT	0.435 411.655 0.485 411.785 ;
		RECT	0.435 411.195 0.485 411.325 ;
		RECT	0.435 413.615 0.485 413.745 ;
		RECT	0.435 250.375 0.485 250.505 ;
		RECT	0.435 249.915 0.485 250.045 ;
		RECT	0.435 252.335 0.485 252.465 ;
		RECT	0.435 253.255 0.485 253.385 ;
		RECT	0.435 252.795 0.485 252.925 ;
		RECT	0.435 255.215 0.485 255.345 ;
		RECT	0.435 256.135 0.485 256.265 ;
		RECT	0.435 255.675 0.485 255.805 ;
		RECT	0.435 258.095 0.485 258.225 ;
		RECT	20.895 186.875 21.075 187.005 ;
		RECT	20.89 221.89 21.02 222.07 ;
		RECT	20.895 227.855 21.075 227.985 ;
		RECT	20.93 192.885 20.98 193.015 ;
		RECT	21.205 188.455 21.385 188.585 ;
		RECT	21.34 190.46 21.39 190.59 ;
		RECT	21.34 193.375 21.39 193.505 ;
		RECT	21.34 194.36 21.39 194.49 ;
		RECT	21.34 196.33 21.39 196.46 ;
		RECT	21.34 197.31 21.39 197.44 ;
		RECT	21.34 198.295 21.39 198.425 ;
		RECT	21.34 201.25 21.39 201.38 ;
		RECT	21.34 208.63 21.39 208.76 ;
		RECT	21.34 209.61 21.39 209.74 ;
		RECT	21.34 213.55 21.39 213.68 ;
		RECT	21.34 216.5 21.39 216.63 ;
		RECT	21.34 217.485 21.39 217.615 ;
		RECT	21.34 218.47 21.39 218.6 ;
		RECT	21.34 220.435 21.39 220.565 ;
		RECT	21.34 221.42 21.39 221.55 ;
		RECT	21.34 224.34 21.39 224.47 ;
		RECT	21.205 226.34 21.385 226.47 ;
		RECT	21.685 187.105 21.865 187.235 ;
		RECT	21.685 227.625 21.865 227.755 ;
		RECT	20.895 187.58 21.075 187.71 ;
		RECT	20.92 227.12 21.05 227.3 ;
		RECT	20.93 189.915 20.98 190.045 ;
		RECT	20.93 193.87 20.98 194 ;
		RECT	20.93 197.805 20.98 197.935 ;
		RECT	20.93 201.74 20.98 201.87 ;
		RECT	20.93 205.675 20.98 205.805 ;
		RECT	20.93 209.12 20.98 209.25 ;
		RECT	20.93 213.055 20.98 213.185 ;
		RECT	20.93 216.995 20.98 217.125 ;
		RECT	20.93 220.93 20.98 221.06 ;
		RECT	20.93 224.88 20.98 225.01 ;
		RECT	15.775 186.875 15.825 187.005 ;
		RECT	20.295 186.875 20.345 187.005 ;
		RECT	15.575 186.875 15.625 187.005 ;
		RECT	20.495 186.875 20.545 187.005 ;
		RECT	15.775 227.855 15.825 227.985 ;
		RECT	20.295 227.855 20.345 227.985 ;
		RECT	15.575 227.855 15.625 227.985 ;
		RECT	20.495 227.855 20.545 227.985 ;
		RECT	21.335 186.645 21.385 186.775 ;
		RECT	21.205 186.645 21.255 186.775 ;
		RECT	21.51 187.105 21.56 187.235 ;
		RECT	21.025 187.965 21.075 188.095 ;
		RECT	20.895 187.965 20.945 188.095 ;
		RECT	21.71 188.74 21.84 188.79 ;
		RECT	21.025 188.945 21.075 189.075 ;
		RECT	20.895 188.945 20.945 189.075 ;
		RECT	21.2 189.44 21.25 189.57 ;
		RECT	21.71 189.72 21.84 189.77 ;
		RECT	21.495 190.19 21.545 190.32 ;
		RECT	21.145 190.19 21.195 190.32 ;
		RECT	20.93 190.915 20.98 191.045 ;
		RECT	21.815 191.41 21.865 191.54 ;
		RECT	21.685 191.41 21.735 191.54 ;
		RECT	20.93 191.9 20.98 192.03 ;
		RECT	20.89 192.185 21.02 192.235 ;
		RECT	21.815 192.39 21.865 192.52 ;
		RECT	21.685 192.39 21.735 192.52 ;
		RECT	20.93 194.855 20.98 194.985 ;
		RECT	21.815 195.345 21.865 195.475 ;
		RECT	21.685 195.345 21.735 195.475 ;
		RECT	20.93 195.835 20.98 195.965 ;
		RECT	20.93 196.82 20.98 196.95 ;
		RECT	20.93 198.79 20.98 198.92 ;
		RECT	21.815 199.28 21.865 199.41 ;
		RECT	21.685 199.28 21.735 199.41 ;
		RECT	20.93 199.77 20.98 199.9 ;
		RECT	21.815 200.265 21.865 200.395 ;
		RECT	21.685 200.265 21.735 200.395 ;
		RECT	20.93 200.755 20.98 200.885 ;
		RECT	21.34 202.235 21.39 202.365 ;
		RECT	20.93 202.73 20.98 202.86 ;
		RECT	21.815 203.215 21.865 203.345 ;
		RECT	21.685 203.215 21.735 203.345 ;
		RECT	20.93 203.71 20.98 203.84 ;
		RECT	21.315 204.185 21.365 204.315 ;
		RECT	21.495 204.495 21.545 204.625 ;
		RECT	21.145 204.495 21.195 204.625 ;
		RECT	21.155 204.81 21.205 204.94 ;
		RECT	21.71 205.47 21.84 205.52 ;
		RECT	21.71 205.965 21.84 206.015 ;
		RECT	20.93 206.66 20.98 206.79 ;
		RECT	21.815 207.15 21.865 207.28 ;
		RECT	21.685 207.15 21.735 207.28 ;
		RECT	21.815 207.645 21.865 207.775 ;
		RECT	21.685 207.645 21.735 207.775 ;
		RECT	20.93 208.135 20.98 208.265 ;
		RECT	21.71 208.915 21.84 208.965 ;
		RECT	21.71 209.405 21.84 209.455 ;
		RECT	21.155 209.925 21.205 210.055 ;
		RECT	21.495 210.27 21.545 210.4 ;
		RECT	21.145 210.27 21.195 210.4 ;
		RECT	20.93 211.085 20.98 211.215 ;
		RECT	21.815 211.58 21.865 211.71 ;
		RECT	21.685 211.58 21.735 211.71 ;
		RECT	20.93 212.075 20.98 212.205 ;
		RECT	21.34 212.565 21.39 212.695 ;
		RECT	20.93 214.04 20.98 214.17 ;
		RECT	21.815 214.535 21.865 214.665 ;
		RECT	21.685 214.535 21.735 214.665 ;
		RECT	20.93 215.025 20.98 215.155 ;
		RECT	21.815 215.515 21.865 215.645 ;
		RECT	21.685 215.515 21.735 215.645 ;
		RECT	20.93 216.01 20.98 216.14 ;
		RECT	20.93 217.975 20.98 218.105 ;
		RECT	20.93 218.96 20.98 219.09 ;
		RECT	21.815 219.455 21.865 219.585 ;
		RECT	21.685 219.455 21.735 219.585 ;
		RECT	20.93 219.945 20.98 220.075 ;
		RECT	20.89 220.72 21.02 220.77 ;
		RECT	20.89 222.2 21.02 222.25 ;
		RECT	21.815 222.405 21.865 222.535 ;
		RECT	21.685 222.405 21.735 222.535 ;
		RECT	20.89 222.69 21.02 222.74 ;
		RECT	20.93 222.895 20.98 223.025 ;
		RECT	21.815 223.355 21.865 223.485 ;
		RECT	21.685 223.355 21.735 223.485 ;
		RECT	20.93 223.88 20.98 224.01 ;
		RECT	21.495 224.61 21.545 224.74 ;
		RECT	21.145 224.61 21.195 224.74 ;
		RECT	21.71 225.155 21.84 225.205 ;
		RECT	21.2 225.355 21.25 225.485 ;
		RECT	21.025 225.85 21.075 225.98 ;
		RECT	20.895 225.85 20.945 225.98 ;
		RECT	21.71 226.135 21.84 226.185 ;
		RECT	21.025 226.835 21.075 226.965 ;
		RECT	20.895 226.835 20.945 226.965 ;
		RECT	21.51 227.625 21.56 227.755 ;
		RECT	21.205 228.085 21.385 228.215 ;
		RECT	15.8 190.915 15.85 191.045 ;
		RECT	15.8 191.9 15.85 192.03 ;
		RECT	15.8 192.185 15.85 192.235 ;
		RECT	15.8 194.855 15.85 194.985 ;
		RECT	15.8 195.835 15.85 195.965 ;
		RECT	15.8 196.82 15.85 196.95 ;
		RECT	15.8 198.79 15.85 198.92 ;
		RECT	15.8 199.77 15.85 199.9 ;
		RECT	15.8 200.755 15.85 200.885 ;
		RECT	15.8 202.73 15.85 202.86 ;
		RECT	15.8 203.71 15.85 203.84 ;
		RECT	15.775 206.66 15.825 206.79 ;
		RECT	15.775 208.135 15.825 208.265 ;
		RECT	15.8 211.085 15.85 211.215 ;
		RECT	15.8 212.075 15.85 212.205 ;
		RECT	15.8 214.04 15.85 214.17 ;
		RECT	15.8 215.025 15.85 215.155 ;
		RECT	15.8 216.01 15.85 216.14 ;
		RECT	15.8 217.975 15.85 218.105 ;
		RECT	15.8 218.96 15.85 219.09 ;
		RECT	15.8 219.945 15.85 220.075 ;
		RECT	15.8 220.72 15.85 220.77 ;
		RECT	15.8 222.895 15.85 223.025 ;
		RECT	15.8 223.88 15.85 224.01 ;
		RECT	20.275 213.03 20.405 213.21 ;
		RECT	20.275 220.905 20.405 221.085 ;
		RECT	20.315 201.74 20.365 201.87 ;
		RECT	20.685 204.185 20.735 204.315 ;
		RECT	20.685 210.61 20.735 210.74 ;
		RECT	20.51 187.965 20.56 188.095 ;
		RECT	20.51 188.945 20.56 189.075 ;
		RECT	20.51 190.915 20.56 191.045 ;
		RECT	20.51 191.9 20.56 192.03 ;
		RECT	20.51 192.185 20.56 192.235 ;
		RECT	20.51 194.855 20.56 194.985 ;
		RECT	20.51 195.835 20.56 195.965 ;
		RECT	20.51 196.82 20.56 196.95 ;
		RECT	20.51 198.79 20.56 198.92 ;
		RECT	20.51 199.77 20.56 199.9 ;
		RECT	20.51 200.755 20.56 200.885 ;
		RECT	20.51 202.73 20.56 202.86 ;
		RECT	20.51 203.71 20.56 203.84 ;
		RECT	20.51 206.66 20.56 206.79 ;
		RECT	20.51 208.135 20.56 208.265 ;
		RECT	20.51 211.085 20.56 211.215 ;
		RECT	20.51 212.075 20.56 212.205 ;
		RECT	20.51 214.04 20.56 214.17 ;
		RECT	20.51 215.025 20.56 215.155 ;
		RECT	20.51 216.01 20.56 216.14 ;
		RECT	20.51 217.975 20.56 218.105 ;
		RECT	20.51 218.96 20.56 219.09 ;
		RECT	20.51 219.945 20.56 220.075 ;
		RECT	20.51 220.72 20.56 220.77 ;
		RECT	20.275 221.89 20.405 222.07 ;
		RECT	20.51 222.895 20.56 223.025 ;
		RECT	20.51 223.88 20.56 224.01 ;
		RECT	20.51 225.85 20.56 225.98 ;
		RECT	20.51 226.835 20.56 226.965 ;
		RECT	15.575 187.965 15.625 188.095 ;
		RECT	15.575 188.945 15.625 189.075 ;
		RECT	15.535 190.915 15.585 191.045 ;
		RECT	15.535 191.9 15.585 192.03 ;
		RECT	15.535 192.185 15.585 192.235 ;
		RECT	15.54 194.855 15.59 194.985 ;
		RECT	15.535 195.835 15.585 195.965 ;
		RECT	15.535 196.82 15.585 196.95 ;
		RECT	15.535 198.79 15.585 198.92 ;
		RECT	15.535 199.77 15.585 199.9 ;
		RECT	15.535 200.755 15.585 200.885 ;
		RECT	15.535 202.73 15.585 202.86 ;
		RECT	15.535 203.71 15.585 203.84 ;
		RECT	15.56 206.66 15.61 206.79 ;
		RECT	15.56 208.135 15.61 208.265 ;
		RECT	15.535 211.085 15.585 211.215 ;
		RECT	15.535 212.075 15.585 212.205 ;
		RECT	15.535 214.04 15.585 214.17 ;
		RECT	15.535 215.025 15.585 215.155 ;
		RECT	15.535 216.01 15.585 216.14 ;
		RECT	15.535 217.975 15.585 218.105 ;
		RECT	15.535 218.96 15.585 219.09 ;
		RECT	15.535 219.945 15.585 220.075 ;
		RECT	15.535 220.72 15.585 220.77 ;
		RECT	15.535 222.895 15.585 223.025 ;
		RECT	15.535 223.88 15.585 224.01 ;
		RECT	15.575 225.85 15.625 225.98 ;
		RECT	15.575 226.835 15.625 226.965 ;
		RECT	15.36 204.185 15.41 204.315 ;
		RECT	15.36 210.61 15.41 210.74 ;
		RECT	15.775 187.965 15.825 188.095 ;
		RECT	16.145 187.965 16.195 188.095 ;
		RECT	16.685 187.965 16.735 188.095 ;
		RECT	17.225 187.965 17.275 188.095 ;
		RECT	17.765 187.965 17.815 188.095 ;
		RECT	18.305 187.965 18.355 188.095 ;
		RECT	18.845 187.965 18.895 188.095 ;
		RECT	19.385 187.965 19.435 188.095 ;
		RECT	19.925 187.965 19.975 188.095 ;
		RECT	15.375 188.74 15.425 188.79 ;
		RECT	15.76 188.945 15.81 189.075 ;
		RECT	16.145 189.44 16.195 189.57 ;
		RECT	16.685 189.44 16.735 189.57 ;
		RECT	17.225 189.44 17.275 189.57 ;
		RECT	17.765 189.44 17.815 189.57 ;
		RECT	18.305 189.44 18.355 189.57 ;
		RECT	18.845 189.44 18.895 189.57 ;
		RECT	19.385 189.44 19.435 189.57 ;
		RECT	19.925 189.44 19.975 189.57 ;
		RECT	15.375 189.72 15.425 189.77 ;
		RECT	15.8 189.915 15.85 190.045 ;
		RECT	15.675 190.19 15.725 190.32 ;
		RECT	16.145 190.19 16.195 190.32 ;
		RECT	16.685 190.19 16.735 190.32 ;
		RECT	17.225 190.19 17.275 190.32 ;
		RECT	17.765 190.19 17.815 190.32 ;
		RECT	18.305 190.19 18.355 190.32 ;
		RECT	18.845 190.19 18.895 190.32 ;
		RECT	19.385 190.19 19.435 190.32 ;
		RECT	19.925 190.19 19.975 190.32 ;
		RECT	15.36 191.41 15.41 191.54 ;
		RECT	15.365 192.39 15.415 192.52 ;
		RECT	15.54 192.885 15.59 193.015 ;
		RECT	15.8 193.87 15.85 194 ;
		RECT	15.365 195.345 15.415 195.475 ;
		RECT	15.8 197.805 15.85 197.935 ;
		RECT	15.36 199.28 15.41 199.41 ;
		RECT	15.36 200.265 15.41 200.395 ;
		RECT	15.8 201.715 15.85 201.765 ;
		RECT	15.8 201.845 15.85 201.895 ;
		RECT	15.36 203.215 15.41 203.345 ;
		RECT	15.675 204.495 15.725 204.625 ;
		RECT	16.145 204.495 16.195 204.625 ;
		RECT	16.685 204.495 16.735 204.625 ;
		RECT	17.225 204.495 17.275 204.625 ;
		RECT	17.765 204.495 17.815 204.625 ;
		RECT	18.305 204.495 18.355 204.625 ;
		RECT	18.845 204.495 18.895 204.625 ;
		RECT	19.385 204.495 19.435 204.625 ;
		RECT	19.925 204.495 19.975 204.625 ;
		RECT	16.145 204.81 16.195 204.94 ;
		RECT	16.685 204.81 16.735 204.94 ;
		RECT	17.225 204.81 17.275 204.94 ;
		RECT	17.765 204.81 17.815 204.94 ;
		RECT	18.305 204.81 18.355 204.94 ;
		RECT	18.845 204.81 18.895 204.94 ;
		RECT	19.385 204.81 19.435 204.94 ;
		RECT	19.925 204.81 19.975 204.94 ;
		RECT	15.375 205.47 15.425 205.52 ;
		RECT	15.775 205.675 15.825 205.805 ;
		RECT	15.375 205.965 15.425 206.015 ;
		RECT	16.145 206.66 16.195 206.79 ;
		RECT	16.685 206.66 16.735 206.79 ;
		RECT	17.225 206.66 17.275 206.79 ;
		RECT	17.765 206.66 17.815 206.79 ;
		RECT	18.305 206.66 18.355 206.79 ;
		RECT	18.845 206.66 18.895 206.79 ;
		RECT	19.385 206.66 19.435 206.79 ;
		RECT	19.925 206.66 19.975 206.79 ;
		RECT	15.365 207.15 15.415 207.28 ;
		RECT	15.365 207.645 15.415 207.775 ;
		RECT	16.145 208.135 16.195 208.265 ;
		RECT	16.685 208.135 16.735 208.265 ;
		RECT	17.225 208.135 17.275 208.265 ;
		RECT	17.765 208.135 17.815 208.265 ;
		RECT	18.305 208.135 18.355 208.265 ;
		RECT	18.845 208.135 18.895 208.265 ;
		RECT	19.385 208.135 19.435 208.265 ;
		RECT	19.925 208.135 19.975 208.265 ;
		RECT	15.375 208.915 15.425 208.965 ;
		RECT	15.775 209.12 15.825 209.25 ;
		RECT	15.375 209.405 15.425 209.455 ;
		RECT	16.145 209.925 16.195 210.055 ;
		RECT	16.685 209.925 16.735 210.055 ;
		RECT	17.225 209.925 17.275 210.055 ;
		RECT	17.765 209.925 17.815 210.055 ;
		RECT	18.305 209.925 18.355 210.055 ;
		RECT	18.845 209.925 18.895 210.055 ;
		RECT	19.385 209.925 19.435 210.055 ;
		RECT	19.925 209.925 19.975 210.055 ;
		RECT	15.675 210.27 15.725 210.4 ;
		RECT	16.145 210.27 16.195 210.4 ;
		RECT	16.685 210.27 16.735 210.4 ;
		RECT	17.225 210.27 17.275 210.4 ;
		RECT	17.765 210.27 17.815 210.4 ;
		RECT	18.305 210.27 18.355 210.4 ;
		RECT	18.845 210.27 18.895 210.4 ;
		RECT	19.385 210.27 19.435 210.4 ;
		RECT	19.925 210.27 19.975 210.4 ;
		RECT	15.36 211.58 15.41 211.71 ;
		RECT	15.8 213.03 15.85 213.08 ;
		RECT	15.8 213.16 15.85 213.21 ;
		RECT	15.365 214.535 15.415 214.665 ;
		RECT	15.365 215.515 15.415 215.645 ;
		RECT	15.8 216.995 15.85 217.125 ;
		RECT	15.365 219.455 15.415 219.585 ;
		RECT	15.8 220.93 15.85 221.06 ;
		RECT	15.54 221.915 15.59 222.045 ;
		RECT	15.375 222.405 15.425 222.535 ;
		RECT	15.36 223.355 15.41 223.485 ;
		RECT	15.675 224.61 15.725 224.74 ;
		RECT	16.145 224.61 16.195 224.74 ;
		RECT	16.685 224.61 16.735 224.74 ;
		RECT	17.225 224.61 17.275 224.74 ;
		RECT	17.765 224.61 17.815 224.74 ;
		RECT	18.305 224.61 18.355 224.74 ;
		RECT	18.845 224.61 18.895 224.74 ;
		RECT	19.385 224.61 19.435 224.74 ;
		RECT	19.925 224.61 19.975 224.74 ;
		RECT	15.8 224.88 15.85 225.01 ;
		RECT	15.375 225.155 15.425 225.205 ;
		RECT	16.145 225.355 16.195 225.485 ;
		RECT	16.685 225.355 16.735 225.485 ;
		RECT	17.225 225.355 17.275 225.485 ;
		RECT	17.765 225.355 17.815 225.485 ;
		RECT	18.305 225.355 18.355 225.485 ;
		RECT	18.845 225.355 18.895 225.485 ;
		RECT	19.385 225.355 19.435 225.485 ;
		RECT	19.925 225.355 19.975 225.485 ;
		RECT	15.76 225.85 15.81 225.98 ;
		RECT	15.375 226.135 15.425 226.185 ;
		RECT	15.76 226.835 15.81 226.965 ;
		RECT	16.145 226.835 16.195 226.965 ;
		RECT	16.685 226.835 16.735 226.965 ;
		RECT	17.225 226.835 17.275 226.965 ;
		RECT	17.765 226.835 17.815 226.965 ;
		RECT	18.305 226.835 18.355 226.965 ;
		RECT	18.845 226.835 18.895 226.965 ;
		RECT	19.385 226.835 19.435 226.965 ;
		RECT	19.925 226.835 19.975 226.965 ;
		RECT	20.275 188.005 20.405 188.055 ;
		RECT	20.66 188.74 20.79 188.79 ;
		RECT	20.695 188.74 20.745 188.79 ;
		RECT	20.3 188.945 20.35 189.075 ;
		RECT	20.66 189.72 20.79 189.77 ;
		RECT	20.275 190.955 20.405 191.005 ;
		RECT	20.695 191.41 20.745 191.54 ;
		RECT	20.275 191.94 20.405 191.99 ;
		RECT	20.275 192.185 20.405 192.235 ;
		RECT	20.695 192.39 20.745 192.52 ;
		RECT	20.51 192.885 20.56 193.015 ;
		RECT	20.275 194.895 20.405 194.945 ;
		RECT	20.695 195.345 20.745 195.475 ;
		RECT	20.275 195.875 20.405 195.925 ;
		RECT	20.275 196.86 20.405 196.91 ;
		RECT	20.275 198.83 20.405 198.88 ;
		RECT	20.695 199.28 20.745 199.41 ;
		RECT	20.275 199.745 20.405 199.795 ;
		RECT	20.275 199.875 20.405 199.925 ;
		RECT	20.695 200.265 20.745 200.395 ;
		RECT	20.275 200.795 20.405 200.845 ;
		RECT	20.275 202.77 20.405 202.82 ;
		RECT	20.695 203.215 20.745 203.345 ;
		RECT	20.275 203.75 20.405 203.8 ;
		RECT	20.66 205.47 20.79 205.52 ;
		RECT	20.695 205.47 20.745 205.52 ;
		RECT	20.66 205.965 20.79 206.015 ;
		RECT	20.695 205.965 20.745 206.015 ;
		RECT	20.275 206.7 20.405 206.75 ;
		RECT	20.695 207.15 20.745 207.28 ;
		RECT	20.695 207.645 20.745 207.775 ;
		RECT	20.275 208.175 20.405 208.225 ;
		RECT	20.66 208.915 20.79 208.965 ;
		RECT	20.695 208.915 20.745 208.965 ;
		RECT	20.66 209.405 20.79 209.455 ;
		RECT	20.695 209.405 20.745 209.455 ;
		RECT	20.275 211.125 20.405 211.175 ;
		RECT	20.695 211.58 20.745 211.71 ;
		RECT	20.275 212.115 20.405 212.165 ;
		RECT	20.275 214.08 20.405 214.13 ;
		RECT	20.695 214.535 20.745 214.665 ;
		RECT	20.275 215 20.405 215.05 ;
		RECT	20.275 215.13 20.405 215.18 ;
		RECT	20.695 215.515 20.745 215.645 ;
		RECT	20.275 216.05 20.405 216.1 ;
		RECT	20.275 218.015 20.405 218.065 ;
		RECT	20.275 219 20.405 219.05 ;
		RECT	20.695 219.455 20.745 219.585 ;
		RECT	20.275 219.985 20.405 220.035 ;
		RECT	20.275 220.72 20.405 220.77 ;
		RECT	20.51 221.915 20.56 222.045 ;
		RECT	20.695 222.405 20.745 222.535 ;
		RECT	20.275 222.87 20.405 222.92 ;
		RECT	20.275 223 20.405 223.05 ;
		RECT	20.695 223.355 20.745 223.485 ;
		RECT	20.275 223.92 20.405 223.97 ;
		RECT	20.66 225.155 20.79 225.205 ;
		RECT	20.695 225.155 20.745 225.205 ;
		RECT	20.275 225.89 20.405 225.94 ;
		RECT	20.695 226.135 20.745 226.185 ;
		RECT	20.275 226.875 20.405 226.925 ;
	END

END rf2_32x128_wm1

END LIBRARY

