



module VX_scheduler (
	input clk,
	input 
	
);

endmodule