`include "VX_raster_define.vh"

module VX_raster_setup #(
    // TODO
) (
    input wire clk,
    input wire reset
    // TODO
);

    // TODO

endmodule