`include "VX_rop_define.vh"

module VX_rop_unit #(  
    parameter CORE_ID = 0
) (
    input wire  clk,
    input wire  reset

    // TODO
);

    // TODO

endmodule