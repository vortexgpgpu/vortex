# Copyright (c) 1993 - 2019 ARM Limited. All Rights Reserved.
# Use of this Software is subject to the terms and conditions of the
# applicable license agreement with ARM Limited.

# PhyVGen V 8.3.0
# ARM Version r4p0
# Creation Date: Sun Oct 20 14:43:11 2019


# Memory Configuration:
# ~~~~~~~~~~~~~~~~~~~~~
#  -activity_factor 50 -atf off -back_biasing off -bits 19 -bmux on
# -bus_notation on -check_instname off -diodes on -drive 6 -ema on -frequency
# 1.0 -instname rf2_256x19_wm0 -left_bus_delim "[" -mux 2 -mvt BASE -name_case
# upper -pipeline off -power_gating off -power_type otc -pwr_gnd_rename
# vddpe:VDDPE,vddce:VDDCE,vsse:VSSE -rcols 2 -redundancy off -retention on
# -right_bus_delim "]" -rrows 0 -ser none -site_def off -top_layer m5-m10
# -words 256 -wp_size 1 -write_mask off -write_thru off -corners
# ff_0p99v_0p99v_125c,ss_0p81v_0p81v_m40c,tt_0p90v_0p90v_25c
# 

VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO rf2_256x19_wm0
	FOREIGN rf2_256x19_wm0 0 0 ;
	SYMMETRY X Y ;
	SIZE 51.405 BY 100.94 ;
	CLASS BLOCK ;
	PIN AA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 32.87 0.25 32.97 ;
			LAYER	M2 ;
			RECT	0 32.87 0.25 32.97 ;
			LAYER	M3 ;
			RECT	0 32.87 0.25 32.97 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[0]

	PIN AA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 35.9 0.25 36 ;
			LAYER	M2 ;
			RECT	0 35.9 0.25 36 ;
			LAYER	M3 ;
			RECT	0 35.9 0.25 36 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[1]

	PIN AA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 37.445 0.25 37.545 ;
			LAYER	M2 ;
			RECT	0 37.445 0.25 37.545 ;
			LAYER	M3 ;
			RECT	0 37.445 0.25 37.545 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[2]

	PIN AA[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 38.93 0.25 39.03 ;
			LAYER	M2 ;
			RECT	0 38.93 0.25 39.03 ;
			LAYER	M3 ;
			RECT	0 38.93 0.25 39.03 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[3]

	PIN AA[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 40.475 0.25 40.575 ;
			LAYER	M2 ;
			RECT	0 40.475 0.25 40.575 ;
			LAYER	M3 ;
			RECT	0 40.475 0.25 40.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[4]

	PIN AA[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 41.96 0.25 42.06 ;
			LAYER	M2 ;
			RECT	0 41.96 0.25 42.06 ;
			LAYER	M3 ;
			RECT	0 41.96 0.25 42.06 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[5]

	PIN AA[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 43.505 0.25 43.605 ;
			LAYER	M2 ;
			RECT	0 43.505 0.25 43.605 ;
			LAYER	M3 ;
			RECT	0 43.505 0.25 43.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[6]

	PIN AA[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 44.99 0.25 45.09 ;
			LAYER	M2 ;
			RECT	0 44.99 0.25 45.09 ;
			LAYER	M3 ;
			RECT	0 44.99 0.25 45.09 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AA[7]

	PIN AB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 65.785 0.25 65.885 ;
			LAYER	M2 ;
			RECT	0 65.785 0.25 65.885 ;
			LAYER	M3 ;
			RECT	0 65.785 0.25 65.885 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[0]

	PIN AB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 62.56 0.25 62.66 ;
			LAYER	M2 ;
			RECT	0 62.56 0.25 62.66 ;
			LAYER	M3 ;
			RECT	0 62.56 0.25 62.66 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[1]

	PIN AB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 61.21 0.25 61.31 ;
			LAYER	M2 ;
			RECT	0 61.21 0.25 61.31 ;
			LAYER	M3 ;
			RECT	0 61.21 0.25 61.31 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[2]

	PIN AB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 59.725 0.25 59.825 ;
			LAYER	M2 ;
			RECT	0 59.725 0.25 59.825 ;
			LAYER	M3 ;
			RECT	0 59.725 0.25 59.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[3]

	PIN AB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 58.18 0.25 58.28 ;
			LAYER	M2 ;
			RECT	0 58.18 0.25 58.28 ;
			LAYER	M3 ;
			RECT	0 58.18 0.25 58.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[4]

	PIN AB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 56.695 0.25 56.795 ;
			LAYER	M2 ;
			RECT	0 56.695 0.25 56.795 ;
			LAYER	M3 ;
			RECT	0 56.695 0.25 56.795 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[5]

	PIN AB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 55.15 0.25 55.25 ;
			LAYER	M2 ;
			RECT	0 55.15 0.25 55.25 ;
			LAYER	M3 ;
			RECT	0 55.15 0.25 55.25 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[6]

	PIN AB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 53.665 0.25 53.765 ;
			LAYER	M2 ;
			RECT	0 53.665 0.25 53.765 ;
			LAYER	M3 ;
			RECT	0 53.665 0.25 53.765 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AB[7]

	PIN AYA[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 33.275 0.25 33.375 ;
			LAYER	M2 ;
			RECT	0 33.275 0.25 33.375 ;
			LAYER	M3 ;
			RECT	0 33.275 0.25 33.375 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[0]

	PIN AYA[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 36.305 0.25 36.405 ;
			LAYER	M2 ;
			RECT	0 36.305 0.25 36.405 ;
			LAYER	M3 ;
			RECT	0 36.305 0.25 36.405 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[1]

	PIN AYA[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 37.04 0.25 37.14 ;
			LAYER	M2 ;
			RECT	0 37.04 0.25 37.14 ;
			LAYER	M3 ;
			RECT	0 37.04 0.25 37.14 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[2]

	PIN AYA[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 39.335 0.25 39.435 ;
			LAYER	M2 ;
			RECT	0 39.335 0.25 39.435 ;
			LAYER	M3 ;
			RECT	0 39.335 0.25 39.435 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[3]

	PIN AYA[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 40.1 0.25 40.2 ;
			LAYER	M2 ;
			RECT	0 40.1 0.25 40.2 ;
			LAYER	M3 ;
			RECT	0 40.1 0.25 40.2 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[4]

	PIN AYA[5]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 42.365 0.25 42.465 ;
			LAYER	M2 ;
			RECT	0 42.365 0.25 42.465 ;
			LAYER	M3 ;
			RECT	0 42.365 0.25 42.465 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[5]

	PIN AYA[6]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 43.305 0.25 43.405 ;
			LAYER	M2 ;
			RECT	0 43.305 0.25 43.405 ;
			LAYER	M3 ;
			RECT	0 43.305 0.25 43.405 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[6]

	PIN AYA[7]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 45.395 0.25 45.495 ;
			LAYER	M2 ;
			RECT	0 45.395 0.25 45.495 ;
			LAYER	M3 ;
			RECT	0 45.395 0.25 45.495 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYA[7]

	PIN AYB[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 65.38 0.25 65.48 ;
			LAYER	M2 ;
			RECT	0 65.38 0.25 65.48 ;
			LAYER	M3 ;
			RECT	0 65.38 0.25 65.48 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[0]

	PIN AYB[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 62.35 0.25 62.45 ;
			LAYER	M2 ;
			RECT	0 62.35 0.25 62.45 ;
			LAYER	M3 ;
			RECT	0 62.35 0.25 62.45 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[1]

	PIN AYB[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 61.585 0.25 61.685 ;
			LAYER	M2 ;
			RECT	0 61.585 0.25 61.685 ;
			LAYER	M3 ;
			RECT	0 61.585 0.25 61.685 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[2]

	PIN AYB[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 59.35 0.25 59.45 ;
			LAYER	M2 ;
			RECT	0 59.35 0.25 59.45 ;
			LAYER	M3 ;
			RECT	0 59.35 0.25 59.45 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[3]

	PIN AYB[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 58.585 0.25 58.685 ;
			LAYER	M2 ;
			RECT	0 58.585 0.25 58.685 ;
			LAYER	M3 ;
			RECT	0 58.585 0.25 58.685 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[4]

	PIN AYB[5]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 56.29 0.25 56.39 ;
			LAYER	M2 ;
			RECT	0 56.29 0.25 56.39 ;
			LAYER	M3 ;
			RECT	0 56.29 0.25 56.39 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[5]

	PIN AYB[6]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 55.525 0.25 55.625 ;
			LAYER	M2 ;
			RECT	0 55.525 0.25 55.625 ;
			LAYER	M3 ;
			RECT	0 55.525 0.25 55.625 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[6]

	PIN AYB[7]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 53.26 0.25 53.36 ;
			LAYER	M2 ;
			RECT	0 53.26 0.25 53.36 ;
			LAYER	M3 ;
			RECT	0 53.26 0.25 53.36 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END AYB[7]

	PIN CENA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 30.11 0.25 30.21 ;
			LAYER	M2 ;
			RECT	0 30.11 0.25 30.21 ;
			LAYER	M3 ;
			RECT	0 30.11 0.25 30.21 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENA

	PIN CENB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 70.305 0.25 70.405 ;
			LAYER	M2 ;
			RECT	0 70.305 0.25 70.405 ;
			LAYER	M3 ;
			RECT	0 70.305 0.25 70.405 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENB

	PIN CENYA
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 28.7 0.25 28.8 ;
			LAYER	M2 ;
			RECT	0 28.7 0.25 28.8 ;
			LAYER	M3 ;
			RECT	0 28.7 0.25 28.8 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENYA

	PIN CENYB
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 70.85 0.25 70.95 ;
			LAYER	M2 ;
			RECT	0 70.85 0.25 70.95 ;
			LAYER	M3 ;
			RECT	0 70.85 0.25 70.95 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CENYB

	PIN CLKA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 39.73 0.25 39.83 ;
			LAYER	M2 ;
			RECT	0 39.73 0.25 39.83 ;
			LAYER	M3 ;
			RECT	0 39.73 0.25 39.83 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CLKA

	PIN CLKB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 60.38 0.25 60.48 ;
			LAYER	M2 ;
			RECT	0 60.38 0.25 60.48 ;
			LAYER	M3 ;
			RECT	0 60.38 0.25 60.48 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END CLKB

	PIN COLLDISN
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 47.9 0.25 48 ;
			LAYER	M2 ;
			RECT	0 47.9 0.25 48 ;
			LAYER	M3 ;
			RECT	0 47.9 0.25 48 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END COLLDISN

	PIN DB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 2.195 0.25 2.295 ;
			LAYER	M2 ;
			RECT	0 2.195 0.25 2.295 ;
			LAYER	M3 ;
			RECT	0 2.195 0.25 2.295 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[0]

	PIN DB[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 75.605 0.25 75.705 ;
			LAYER	M2 ;
			RECT	0 75.605 0.25 75.705 ;
			LAYER	M3 ;
			RECT	0 75.605 0.25 75.705 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[10]

	PIN DB[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 78.485 0.25 78.585 ;
			LAYER	M2 ;
			RECT	0 78.485 0.25 78.585 ;
			LAYER	M3 ;
			RECT	0 78.485 0.25 78.585 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[11]

	PIN DB[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 81.365 0.25 81.465 ;
			LAYER	M2 ;
			RECT	0 81.365 0.25 81.465 ;
			LAYER	M3 ;
			RECT	0 81.365 0.25 81.465 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[12]

	PIN DB[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 84.245 0.25 84.345 ;
			LAYER	M2 ;
			RECT	0 84.245 0.25 84.345 ;
			LAYER	M3 ;
			RECT	0 84.245 0.25 84.345 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[13]

	PIN DB[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 87.125 0.25 87.225 ;
			LAYER	M2 ;
			RECT	0 87.125 0.25 87.225 ;
			LAYER	M3 ;
			RECT	0 87.125 0.25 87.225 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[14]

	PIN DB[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 90.005 0.25 90.105 ;
			LAYER	M2 ;
			RECT	0 90.005 0.25 90.105 ;
			LAYER	M3 ;
			RECT	0 90.005 0.25 90.105 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[15]

	PIN DB[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 92.885 0.25 92.985 ;
			LAYER	M2 ;
			RECT	0 92.885 0.25 92.985 ;
			LAYER	M3 ;
			RECT	0 92.885 0.25 92.985 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[16]

	PIN DB[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 95.765 0.25 95.865 ;
			LAYER	M2 ;
			RECT	0 95.765 0.25 95.865 ;
			LAYER	M3 ;
			RECT	0 95.765 0.25 95.865 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[17]

	PIN DB[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 98.645 0.25 98.745 ;
			LAYER	M2 ;
			RECT	0 98.645 0.25 98.745 ;
			LAYER	M3 ;
			RECT	0 98.645 0.25 98.745 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[18]

	PIN DB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 5.075 0.25 5.175 ;
			LAYER	M2 ;
			RECT	0 5.075 0.25 5.175 ;
			LAYER	M3 ;
			RECT	0 5.075 0.25 5.175 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[1]

	PIN DB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 7.955 0.25 8.055 ;
			LAYER	M2 ;
			RECT	0 7.955 0.25 8.055 ;
			LAYER	M3 ;
			RECT	0 7.955 0.25 8.055 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[2]

	PIN DB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 10.835 0.25 10.935 ;
			LAYER	M2 ;
			RECT	0 10.835 0.25 10.935 ;
			LAYER	M3 ;
			RECT	0 10.835 0.25 10.935 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[3]

	PIN DB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 13.715 0.25 13.815 ;
			LAYER	M2 ;
			RECT	0 13.715 0.25 13.815 ;
			LAYER	M3 ;
			RECT	0 13.715 0.25 13.815 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[4]

	PIN DB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 16.595 0.25 16.695 ;
			LAYER	M2 ;
			RECT	0 16.595 0.25 16.695 ;
			LAYER	M3 ;
			RECT	0 16.595 0.25 16.695 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[5]

	PIN DB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 19.475 0.25 19.575 ;
			LAYER	M2 ;
			RECT	0 19.475 0.25 19.575 ;
			LAYER	M3 ;
			RECT	0 19.475 0.25 19.575 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[6]

	PIN DB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 22.355 0.25 22.455 ;
			LAYER	M2 ;
			RECT	0 22.355 0.25 22.455 ;
			LAYER	M3 ;
			RECT	0 22.355 0.25 22.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[7]

	PIN DB[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 25.235 0.25 25.335 ;
			LAYER	M2 ;
			RECT	0 25.235 0.25 25.335 ;
			LAYER	M3 ;
			RECT	0 25.235 0.25 25.335 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[8]

	PIN DB[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 72.725 0.25 72.825 ;
			LAYER	M2 ;
			RECT	0 72.725 0.25 72.825 ;
			LAYER	M3 ;
			RECT	0 72.725 0.25 72.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DB[9]

	PIN DFTRAMBYP
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 67.3 0.25 67.4 ;
			LAYER	M2 ;
			RECT	0 67.3 0.25 67.4 ;
			LAYER	M3 ;
			RECT	0 67.3 0.25 67.4 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END DFTRAMBYP

	PIN EMAA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 41.37 0.25 41.47 ;
			LAYER	M2 ;
			RECT	0 41.37 0.25 41.47 ;
			LAYER	M3 ;
			RECT	0 41.37 0.25 41.47 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAA[0]

	PIN EMAA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 41.17 0.25 41.27 ;
			LAYER	M2 ;
			RECT	0 41.17 0.25 41.27 ;
			LAYER	M3 ;
			RECT	0 41.17 0.25 41.27 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAA[1]

	PIN EMAA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 43.105 0.25 43.205 ;
			LAYER	M2 ;
			RECT	0 43.105 0.25 43.205 ;
			LAYER	M3 ;
			RECT	0 43.105 0.25 43.205 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAA[2]

	PIN EMAB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 55.905 0.25 56.005 ;
			LAYER	M2 ;
			RECT	0 55.905 0.25 56.005 ;
			LAYER	M3 ;
			RECT	0 55.905 0.25 56.005 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAB[0]

	PIN EMAB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 56.905 0.25 57.005 ;
			LAYER	M2 ;
			RECT	0 56.905 0.25 57.005 ;
			LAYER	M3 ;
			RECT	0 56.905 0.25 57.005 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAB[1]

	PIN EMAB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 54.425 0.25 54.525 ;
			LAYER	M2 ;
			RECT	0 54.425 0.25 54.525 ;
			LAYER	M3 ;
			RECT	0 54.425 0.25 54.525 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMAB[2]

	PIN EMASA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 29.05 0.25 29.15 ;
			LAYER	M2 ;
			RECT	0 29.05 0.25 29.15 ;
			LAYER	M3 ;
			RECT	0 29.05 0.25 29.15 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END EMASA

	PIN QA[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 2.455 0.25 2.555 ;
			LAYER	M2 ;
			RECT	0 2.455 0.25 2.555 ;
			LAYER	M3 ;
			RECT	0 2.455 0.25 2.555 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[0]

	PIN QA[10]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 75.345 0.25 75.445 ;
			LAYER	M2 ;
			RECT	0 75.345 0.25 75.445 ;
			LAYER	M3 ;
			RECT	0 75.345 0.25 75.445 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[10]

	PIN QA[11]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 78.225 0.25 78.325 ;
			LAYER	M2 ;
			RECT	0 78.225 0.25 78.325 ;
			LAYER	M3 ;
			RECT	0 78.225 0.25 78.325 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[11]

	PIN QA[12]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 81.105 0.25 81.205 ;
			LAYER	M2 ;
			RECT	0 81.105 0.25 81.205 ;
			LAYER	M3 ;
			RECT	0 81.105 0.25 81.205 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[12]

	PIN QA[13]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 83.985 0.25 84.085 ;
			LAYER	M2 ;
			RECT	0 83.985 0.25 84.085 ;
			LAYER	M3 ;
			RECT	0 83.985 0.25 84.085 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[13]

	PIN QA[14]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 86.865 0.25 86.965 ;
			LAYER	M2 ;
			RECT	0 86.865 0.25 86.965 ;
			LAYER	M3 ;
			RECT	0 86.865 0.25 86.965 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[14]

	PIN QA[15]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 89.745 0.25 89.845 ;
			LAYER	M2 ;
			RECT	0 89.745 0.25 89.845 ;
			LAYER	M3 ;
			RECT	0 89.745 0.25 89.845 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[15]

	PIN QA[16]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 92.625 0.25 92.725 ;
			LAYER	M2 ;
			RECT	0 92.625 0.25 92.725 ;
			LAYER	M3 ;
			RECT	0 92.625 0.25 92.725 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[16]

	PIN QA[17]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 95.505 0.25 95.605 ;
			LAYER	M2 ;
			RECT	0 95.505 0.25 95.605 ;
			LAYER	M3 ;
			RECT	0 95.505 0.25 95.605 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[17]

	PIN QA[18]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 98.385 0.25 98.485 ;
			LAYER	M2 ;
			RECT	0 98.385 0.25 98.485 ;
			LAYER	M3 ;
			RECT	0 98.385 0.25 98.485 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[18]

	PIN QA[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 5.335 0.25 5.435 ;
			LAYER	M2 ;
			RECT	0 5.335 0.25 5.435 ;
			LAYER	M3 ;
			RECT	0 5.335 0.25 5.435 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[1]

	PIN QA[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 8.215 0.25 8.315 ;
			LAYER	M2 ;
			RECT	0 8.215 0.25 8.315 ;
			LAYER	M3 ;
			RECT	0 8.215 0.25 8.315 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[2]

	PIN QA[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 11.095 0.25 11.195 ;
			LAYER	M2 ;
			RECT	0 11.095 0.25 11.195 ;
			LAYER	M3 ;
			RECT	0 11.095 0.25 11.195 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[3]

	PIN QA[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 13.975 0.25 14.075 ;
			LAYER	M2 ;
			RECT	0 13.975 0.25 14.075 ;
			LAYER	M3 ;
			RECT	0 13.975 0.25 14.075 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[4]

	PIN QA[5]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 16.855 0.25 16.955 ;
			LAYER	M2 ;
			RECT	0 16.855 0.25 16.955 ;
			LAYER	M3 ;
			RECT	0 16.855 0.25 16.955 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[5]

	PIN QA[6]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 19.735 0.25 19.835 ;
			LAYER	M2 ;
			RECT	0 19.735 0.25 19.835 ;
			LAYER	M3 ;
			RECT	0 19.735 0.25 19.835 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[6]

	PIN QA[7]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 22.615 0.25 22.715 ;
			LAYER	M2 ;
			RECT	0 22.615 0.25 22.715 ;
			LAYER	M3 ;
			RECT	0 22.615 0.25 22.715 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[7]

	PIN QA[8]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 25.495 0.25 25.595 ;
			LAYER	M2 ;
			RECT	0 25.495 0.25 25.595 ;
			LAYER	M3 ;
			RECT	0 25.495 0.25 25.595 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[8]

	PIN QA[9]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 72.465 0.25 72.565 ;
			LAYER	M2 ;
			RECT	0 72.465 0.25 72.565 ;
			LAYER	M3 ;
			RECT	0 72.465 0.25 72.565 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END QA[9]

	PIN RET1N
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 29.71 0.25 29.81 ;
			LAYER	M2 ;
			RECT	0 29.71 0.25 29.81 ;
			LAYER	M3 ;
			RECT	0 29.71 0.25 29.81 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END RET1N

	PIN SEA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 47.5 0.25 47.6 ;
			LAYER	M2 ;
			RECT	0 47.5 0.25 47.6 ;
			LAYER	M3 ;
			RECT	0 47.5 0.25 47.6 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SEA

	PIN SEB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 50.335 0.25 50.435 ;
			LAYER	M2 ;
			RECT	0 50.335 0.25 50.435 ;
			LAYER	M3 ;
			RECT	0 50.335 0.25 50.435 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SEB

	PIN SIA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 47.7 0.25 47.8 ;
			LAYER	M2 ;
			RECT	0 47.7 0.25 47.8 ;
			LAYER	M3 ;
			RECT	0 47.7 0.25 47.8 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIA[0]

	PIN SIA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 48.67 0.25 48.77 ;
			LAYER	M2 ;
			RECT	0 48.67 0.25 48.77 ;
			LAYER	M3 ;
			RECT	0 48.67 0.25 48.77 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIA[1]

	PIN SIB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 44.275 0.25 44.375 ;
			LAYER	M2 ;
			RECT	0 44.275 0.25 44.375 ;
			LAYER	M3 ;
			RECT	0 44.275 0.25 44.375 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIB[0]

	PIN SIB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 61.925 0.25 62.025 ;
			LAYER	M2 ;
			RECT	0 61.925 0.25 62.025 ;
			LAYER	M3 ;
			RECT	0 61.925 0.25 62.025 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SIB[1]

	PIN SOA[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 0.36 0.25 0.46 ;
			LAYER	M2 ;
			RECT	0 0.36 0.25 0.46 ;
			LAYER	M3 ;
			RECT	0 0.36 0.25 0.46 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOA[0]

	PIN SOA[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 100.48 0.25 100.58 ;
			LAYER	M2 ;
			RECT	0 100.48 0.25 100.58 ;
			LAYER	M3 ;
			RECT	0 100.48 0.25 100.58 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOA[1]

	PIN SOB[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 0.09 0.25 0.19 ;
			LAYER	M2 ;
			RECT	0 0.09 0.25 0.19 ;
			LAYER	M3 ;
			RECT	0 0.09 0.25 0.19 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOB[0]

	PIN SOB[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 100.75 0.25 100.85 ;
			LAYER	M2 ;
			RECT	0 100.75 0.25 100.85 ;
			LAYER	M3 ;
			RECT	0 100.75 0.25 100.85 ;
		END

		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END SOB[1]

	PIN TAA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 32.355 0.25 32.455 ;
			LAYER	M2 ;
			RECT	0 32.355 0.25 32.455 ;
			LAYER	M3 ;
			RECT	0 32.355 0.25 32.455 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[0]

	PIN TAA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 35.385 0.25 35.485 ;
			LAYER	M2 ;
			RECT	0 35.385 0.25 35.485 ;
			LAYER	M3 ;
			RECT	0 35.385 0.25 35.485 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[1]

	PIN TAA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 37.96 0.25 38.06 ;
			LAYER	M2 ;
			RECT	0 37.96 0.25 38.06 ;
			LAYER	M3 ;
			RECT	0 37.96 0.25 38.06 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[2]

	PIN TAA[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 38.445 0.25 38.545 ;
			LAYER	M2 ;
			RECT	0 38.445 0.25 38.545 ;
			LAYER	M3 ;
			RECT	0 38.445 0.25 38.545 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[3]

	PIN TAA[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 40.96 0.25 41.06 ;
			LAYER	M2 ;
			RECT	0 40.96 0.25 41.06 ;
			LAYER	M3 ;
			RECT	0 40.96 0.25 41.06 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[4]

	PIN TAA[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 41.57 0.25 41.67 ;
			LAYER	M2 ;
			RECT	0 41.57 0.25 41.67 ;
			LAYER	M3 ;
			RECT	0 41.57 0.25 41.67 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[5]

	PIN TAA[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 43.99 0.25 44.09 ;
			LAYER	M2 ;
			RECT	0 43.99 0.25 44.09 ;
			LAYER	M3 ;
			RECT	0 43.99 0.25 44.09 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[6]

	PIN TAA[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 44.505 0.25 44.605 ;
			LAYER	M2 ;
			RECT	0 44.505 0.25 44.605 ;
			LAYER	M3 ;
			RECT	0 44.505 0.25 44.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAA[7]

	PIN TAB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 66.27 0.25 66.37 ;
			LAYER	M2 ;
			RECT	0 66.27 0.25 66.37 ;
			LAYER	M3 ;
			RECT	0 66.27 0.25 66.37 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[0]

	PIN TAB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 63.24 0.25 63.34 ;
			LAYER	M2 ;
			RECT	0 63.24 0.25 63.34 ;
			LAYER	M3 ;
			RECT	0 63.24 0.25 63.34 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[1]

	PIN TAB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 60.725 0.25 60.825 ;
			LAYER	M2 ;
			RECT	0 60.725 0.25 60.825 ;
			LAYER	M3 ;
			RECT	0 60.725 0.25 60.825 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[2]

	PIN TAB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 60.18 0.25 60.28 ;
			LAYER	M2 ;
			RECT	0 60.18 0.25 60.28 ;
			LAYER	M3 ;
			RECT	0 60.18 0.25 60.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[3]

	PIN TAB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 57.695 0.25 57.795 ;
			LAYER	M2 ;
			RECT	0 57.695 0.25 57.795 ;
			LAYER	M3 ;
			RECT	0 57.695 0.25 57.795 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[4]

	PIN TAB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 57.18 0.25 57.28 ;
			LAYER	M2 ;
			RECT	0 57.18 0.25 57.28 ;
			LAYER	M3 ;
			RECT	0 57.18 0.25 57.28 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[5]

	PIN TAB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 54.66 0.25 54.76 ;
			LAYER	M2 ;
			RECT	0 54.66 0.25 54.76 ;
			LAYER	M3 ;
			RECT	0 54.66 0.25 54.76 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[6]

	PIN TAB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 54.15 0.25 54.25 ;
			LAYER	M2 ;
			RECT	0 54.15 0.25 54.25 ;
			LAYER	M3 ;
			RECT	0 54.15 0.25 54.25 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TAB[7]

	PIN TCENA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 29.91 0.25 30.01 ;
			LAYER	M2 ;
			RECT	0 29.91 0.25 30.01 ;
			LAYER	M3 ;
			RECT	0 29.91 0.25 30.01 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TCENA

	PIN TCENB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 69.91 0.25 70.01 ;
			LAYER	M2 ;
			RECT	0 69.91 0.25 70.01 ;
			LAYER	M3 ;
			RECT	0 69.91 0.25 70.01 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TCENB

	PIN TDB[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 1.465 0.25 1.565 ;
			LAYER	M2 ;
			RECT	0 1.465 0.25 1.565 ;
			LAYER	M3 ;
			RECT	0 1.465 0.25 1.565 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[0]

	PIN TDB[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 76.335 0.25 76.435 ;
			LAYER	M2 ;
			RECT	0 76.335 0.25 76.435 ;
			LAYER	M3 ;
			RECT	0 76.335 0.25 76.435 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[10]

	PIN TDB[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 79.215 0.25 79.315 ;
			LAYER	M2 ;
			RECT	0 79.215 0.25 79.315 ;
			LAYER	M3 ;
			RECT	0 79.215 0.25 79.315 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[11]

	PIN TDB[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 82.095 0.25 82.195 ;
			LAYER	M2 ;
			RECT	0 82.095 0.25 82.195 ;
			LAYER	M3 ;
			RECT	0 82.095 0.25 82.195 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[12]

	PIN TDB[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 84.975 0.25 85.075 ;
			LAYER	M2 ;
			RECT	0 84.975 0.25 85.075 ;
			LAYER	M3 ;
			RECT	0 84.975 0.25 85.075 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[13]

	PIN TDB[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 87.855 0.25 87.955 ;
			LAYER	M2 ;
			RECT	0 87.855 0.25 87.955 ;
			LAYER	M3 ;
			RECT	0 87.855 0.25 87.955 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[14]

	PIN TDB[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 90.735 0.25 90.835 ;
			LAYER	M2 ;
			RECT	0 90.735 0.25 90.835 ;
			LAYER	M3 ;
			RECT	0 90.735 0.25 90.835 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[15]

	PIN TDB[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 93.615 0.25 93.715 ;
			LAYER	M2 ;
			RECT	0 93.615 0.25 93.715 ;
			LAYER	M3 ;
			RECT	0 93.615 0.25 93.715 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[16]

	PIN TDB[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 96.495 0.25 96.595 ;
			LAYER	M2 ;
			RECT	0 96.495 0.25 96.595 ;
			LAYER	M3 ;
			RECT	0 96.495 0.25 96.595 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[17]

	PIN TDB[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 99.375 0.25 99.475 ;
			LAYER	M2 ;
			RECT	0 99.375 0.25 99.475 ;
			LAYER	M3 ;
			RECT	0 99.375 0.25 99.475 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[18]

	PIN TDB[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 4.345 0.25 4.445 ;
			LAYER	M2 ;
			RECT	0 4.345 0.25 4.445 ;
			LAYER	M3 ;
			RECT	0 4.345 0.25 4.445 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[1]

	PIN TDB[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 7.225 0.25 7.325 ;
			LAYER	M2 ;
			RECT	0 7.225 0.25 7.325 ;
			LAYER	M3 ;
			RECT	0 7.225 0.25 7.325 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[2]

	PIN TDB[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 10.105 0.25 10.205 ;
			LAYER	M2 ;
			RECT	0 10.105 0.25 10.205 ;
			LAYER	M3 ;
			RECT	0 10.105 0.25 10.205 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[3]

	PIN TDB[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 12.985 0.25 13.085 ;
			LAYER	M2 ;
			RECT	0 12.985 0.25 13.085 ;
			LAYER	M3 ;
			RECT	0 12.985 0.25 13.085 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[4]

	PIN TDB[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 15.865 0.25 15.965 ;
			LAYER	M2 ;
			RECT	0 15.865 0.25 15.965 ;
			LAYER	M3 ;
			RECT	0 15.865 0.25 15.965 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[5]

	PIN TDB[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 18.745 0.25 18.845 ;
			LAYER	M2 ;
			RECT	0 18.745 0.25 18.845 ;
			LAYER	M3 ;
			RECT	0 18.745 0.25 18.845 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[6]

	PIN TDB[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 21.625 0.25 21.725 ;
			LAYER	M2 ;
			RECT	0 21.625 0.25 21.725 ;
			LAYER	M3 ;
			RECT	0 21.625 0.25 21.725 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[7]

	PIN TDB[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 24.505 0.25 24.605 ;
			LAYER	M2 ;
			RECT	0 24.505 0.25 24.605 ;
			LAYER	M3 ;
			RECT	0 24.505 0.25 24.605 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[8]

	PIN TDB[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 73.455 0.25 73.555 ;
			LAYER	M2 ;
			RECT	0 73.455 0.25 73.555 ;
			LAYER	M3 ;
			RECT	0 73.455 0.25 73.555 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TDB[9]

	PIN TENA
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 32.05 0.25 32.15 ;
			LAYER	M2 ;
			RECT	0 32.05 0.25 32.15 ;
			LAYER	M3 ;
			RECT	0 32.05 0.25 32.15 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TENA

	PIN TENB
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	M1 ;
			RECT	0 66.525 0.25 66.625 ;
			LAYER	M2 ;
			RECT	0 66.525 0.25 66.625 ;
			LAYER	M3 ;
			RECT	0 66.525 0.25 66.625 ;
		END

		ANTENNAGATEAREA 0.014 ;
		ANTENNADIFFAREA 0.018 ;
		ANTENNAPARTIALMETALAREA 0.025 ;
	END TENB

	PIN VDDCE
		USE POWER ;
		DIRECTION INOUT ;
		PORT
			LAYER	M4 ;
			RECT	0 26.335 51.405 26.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 23.455 51.405 23.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 20.575 51.405 20.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 17.695 51.405 17.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 97.495 51.405 97.645 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 94.615 51.405 94.765 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 91.735 51.405 91.885 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 88.855 51.405 89.005 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 85.975 51.405 86.125 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 83.095 51.405 83.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 80.215 51.405 80.365 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 77.335 51.405 77.485 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 74.455 51.405 74.605 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 71.575 51.405 71.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 14.815 51.405 14.965 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 11.935 51.405 12.085 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.055 51.405 9.205 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.175 51.405 6.325 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.295 51.405 3.445 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 48.72 51.405 48.91 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 49.215 51.405 49.405 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 53.15 51.405 53.34 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 56.105 51.405 56.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 57.085 51.405 57.275 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 61.025 51.405 61.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 63.975 51.405 64.165 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 64.925 51.405 65.115 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.98 51.405 33.17 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 33.96 51.405 34.15 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 36.915 51.405 37.105 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 40.85 51.405 41.04 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 41.835 51.405 42.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 44.785 51.405 44.975 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 100.375 51.405 100.525 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.415 51.405 0.565 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 28.695 51.405 28.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 69.215 51.405 69.365 ;
		END

	END VDDCE

	PIN VDDPE
		USE POWER ;
		DIRECTION INOUT ;
		PORT
			LAYER	M4 ;
			RECT	0 30.025 51.405 30.215 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.03 51.405 32.22 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 34.945 51.405 35.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 35.93 51.405 36.12 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 37.9 51.405 38.09 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 38.88 51.405 39.07 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 39.865 51.405 40.055 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 42.82 51.405 43.01 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 23.915 51.405 24.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 21.035 51.405 21.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 18.155 51.405 18.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 99.915 51.405 100.065 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 97.035 51.405 97.185 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 94.155 51.405 94.305 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 91.275 51.405 91.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 88.395 51.405 88.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 85.515 51.405 85.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 82.635 51.405 82.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 79.755 51.405 79.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 76.875 51.405 77.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 73.995 51.405 74.145 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 15.275 51.405 15.425 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 12.395 51.405 12.545 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.515 51.405 9.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.635 51.405 6.785 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.755 51.405 3.905 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.875 51.405 1.025 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 46.755 51.405 46.945 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 47.74 51.405 47.93 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 50.2 51.405 50.39 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 51.18 51.405 51.37 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 55.12 51.405 55.31 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 58.07 51.405 58.26 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 59.055 51.405 59.245 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 60.04 51.405 60.23 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 62.005 51.405 62.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 62.99 51.405 63.18 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 65.91 51.405 66.1 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 67.91 51.405 68.1 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 100.605 51.405 100.755 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.185 51.405 0.335 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 28.235 51.405 28.385 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 69.675 51.405 69.825 ;
		END

	END VDDPE

	PIN VSSE
		USE GROUND ;
		DIRECTION INOUT ;
		PORT
			LAYER	M4 ;
			RECT	0 100.145 51.405 100.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 0.645 51.405 0.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 28.465 51.405 28.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 69.445 51.405 69.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 97.265 51.405 97.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 94.385 51.405 94.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 26.565 51.405 26.715 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 23.685 51.405 23.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 20.805 51.405 20.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 17.925 51.405 18.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 15.045 51.405 15.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 12.165 51.405 12.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.285 51.405 9.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.405 51.405 6.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 91.505 51.405 91.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.525 51.405 3.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 88.625 51.405 88.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 85.745 51.405 85.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 82.865 51.405 83.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 79.985 51.405 80.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 77.105 51.405 77.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 74.225 51.405 74.375 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 71.345 51.405 71.495 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 99.685 51.405 99.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 24.145 51.405 24.295 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 21.265 51.405 21.415 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 18.385 51.405 18.535 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 93.925 51.405 94.075 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 15.505 51.405 15.655 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 12.625 51.405 12.775 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 9.745 51.405 9.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 6.865 51.405 7.015 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 3.985 51.405 4.135 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 1.105 51.405 1.255 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 91.045 51.405 91.195 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 88.165 51.405 88.315 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 85.285 51.405 85.435 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 82.405 51.405 82.555 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 79.525 51.405 79.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 76.645 51.405 76.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 73.765 51.405 73.915 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 96.805 51.405 96.955 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 29.535 51.405 29.725 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 30.515 51.405 30.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 32.485 51.405 32.675 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 33.47 51.405 33.66 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 36.425 51.405 36.615 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 37.405 51.405 37.595 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 38.39 51.405 38.58 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 40.36 51.405 40.55 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 41.33 51.405 41.54 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 42.325 51.405 42.515 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 44.3 51.405 44.49 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 45.28 51.405 45.47 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 48.23 51.405 48.42 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 49.705 51.405 49.895 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 52.655 51.405 52.845 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 53.645 51.405 53.835 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 55.61 51.405 55.8 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 56.585 51.405 56.795 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 57.58 51.405 57.77 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 59.545 51.405 59.735 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 60.53 51.405 60.72 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 61.515 51.405 61.705 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 64.455 51.405 64.665 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 65.45 51.405 65.64 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 67.42 51.405 67.61 ;
		END

		PORT
			LAYER	M4 ;
			RECT	0 68.405 51.405 68.595 ;
		END

	END VSSE

	OBS
		LAYER	M1 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0.35 51.085 100.59 ;
		RECT	0 0.56 0.32 1.365 ;
		RECT	0 1.665 0.32 2.095 ;
		RECT	0 2.655 0.32 4.245 ;
		RECT	0 4.545 0.32 4.975 ;
		RECT	0 5.535 0.32 7.125 ;
		RECT	0 7.425 0.32 7.855 ;
		RECT	0 8.415 0.32 10.005 ;
		RECT	0 10.305 0.32 10.735 ;
		RECT	0 11.295 0.32 12.885 ;
		RECT	0 13.185 0.32 13.615 ;
		RECT	0 14.175 0.32 15.765 ;
		RECT	0 16.065 0.32 16.495 ;
		RECT	0 17.055 0.32 18.645 ;
		RECT	0 18.945 0.32 19.375 ;
		RECT	0 19.935 0.32 21.525 ;
		RECT	0 21.825 0.32 22.255 ;
		RECT	0 22.815 0.32 24.405 ;
		RECT	0 24.705 0.32 25.135 ;
		RECT	0 25.695 0.32 28.6 ;
		RECT	0 28.9 0.32 28.95 ;
		RECT	0 29.25 0.32 29.61 ;
		RECT	0 30.31 0.32 31.95 ;
		RECT	0 32.555 0.32 32.77 ;
		RECT	0 33.07 0.32 33.175 ;
		RECT	0 33.475 0.32 35.285 ;
		RECT	0 35.585 0.32 35.8 ;
		RECT	0 36.1 0.32 36.205 ;
		RECT	0 36.505 0.32 36.94 ;
		RECT	0 37.24 0.32 37.345 ;
		RECT	0 37.645 0.32 37.86 ;
		RECT	0 38.16 0.32 38.345 ;
		RECT	0 38.645 0.32 38.83 ;
		RECT	0 39.13 0.32 39.235 ;
		RECT	0 39.535 0.32 39.63 ;
		RECT	0 39.93 0.32 40 ;
		RECT	0 40.3 0.32 40.375 ;
		RECT	0 40.675 0.32 40.86 ;
		RECT	0 41.77 0.32 41.86 ;
		RECT	0 42.16 0.32 42.265 ;
		RECT	0 42.565 0.32 43.005 ;
		RECT	0 43.705 0.32 43.89 ;
		RECT	0 44.705 0.32 44.89 ;
		RECT	0 45.19 0.32 45.295 ;
		RECT	0 45.595 0.32 47.4 ;
		RECT	0 48.1 0.32 48.57 ;
		RECT	0 48.87 0.32 50.235 ;
		RECT	0 50.535 0.32 53.16 ;
		RECT	0 53.46 0.32 53.565 ;
		RECT	0 53.865 0.32 54.05 ;
		RECT	0 54.86 0.32 55.05 ;
		RECT	0 55.35 0.32 55.425 ;
		RECT	0 55.725 0.32 55.805 ;
		RECT	0 56.105 0.32 56.19 ;
		RECT	0 56.49 0.32 56.595 ;
		RECT	0 57.38 0.32 57.595 ;
		RECT	0 57.895 0.32 58.08 ;
		RECT	0 58.38 0.32 58.485 ;
		RECT	0 58.785 0.32 59.25 ;
		RECT	0 59.55 0.32 59.625 ;
		RECT	0 59.925 0.32 60.08 ;
		RECT	0 60.925 0.32 61.11 ;
		RECT	0 61.41 0.32 61.485 ;
		RECT	0 62.125 0.32 62.25 ;
		RECT	0 62.76 0.32 63.14 ;
		RECT	0 63.44 0.32 65.28 ;
		RECT	0 65.58 0.32 65.685 ;
		RECT	0 65.985 0.32 66.17 ;
		RECT	0 66.725 0.32 67.2 ;
		RECT	0 67.5 0.32 69.81 ;
		RECT	0 70.11 0.32 70.205 ;
		RECT	0 70.505 0.32 70.75 ;
		RECT	0 71.05 0.32 72.365 ;
		RECT	0 72.925 0.32 73.355 ;
		RECT	0 73.655 0.32 75.245 ;
		RECT	0 75.805 0.32 76.235 ;
		RECT	0 76.535 0.32 78.125 ;
		RECT	0 78.685 0.32 79.115 ;
		RECT	0 79.415 0.32 81.005 ;
		RECT	0 81.565 0.32 81.995 ;
		RECT	0 82.295 0.32 83.885 ;
		RECT	0 84.445 0.32 84.875 ;
		RECT	0 85.175 0.32 86.765 ;
		RECT	0 87.325 0.32 87.755 ;
		RECT	0 88.055 0.32 89.645 ;
		RECT	0 90.205 0.32 90.635 ;
		RECT	0 90.935 0.32 92.525 ;
		RECT	0 93.085 0.32 93.515 ;
		RECT	0 93.815 0.32 95.405 ;
		RECT	0 95.965 0.32 96.395 ;
		RECT	0 96.695 0.32 98.285 ;
		RECT	0 98.845 0.32 99.275 ;
		RECT	0 99.575 0.32 100.38 ;
		RECT	51.085 0 51.405 100.94 ;
		RECT	0.32 0 51.085 0.35 ;
		RECT	0.32 100.59 51.085 100.94 ;
		LAYER	M2 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0.35 51.085 100.59 ;
		RECT	0 0.56 0.32 1.365 ;
		RECT	0 1.665 0.32 2.095 ;
		RECT	0 2.655 0.32 4.245 ;
		RECT	0 4.545 0.32 4.975 ;
		RECT	0 5.535 0.32 7.125 ;
		RECT	0 7.425 0.32 7.855 ;
		RECT	0 8.415 0.32 10.005 ;
		RECT	0 10.305 0.32 10.735 ;
		RECT	0 11.295 0.32 12.885 ;
		RECT	0 13.185 0.32 13.615 ;
		RECT	0 14.175 0.32 15.765 ;
		RECT	0 16.065 0.32 16.495 ;
		RECT	0 17.055 0.32 18.645 ;
		RECT	0 18.945 0.32 19.375 ;
		RECT	0 19.935 0.32 21.525 ;
		RECT	0 21.825 0.32 22.255 ;
		RECT	0 22.815 0.32 24.405 ;
		RECT	0 24.705 0.32 25.135 ;
		RECT	0 25.695 0.32 28.6 ;
		RECT	0 28.9 0.32 28.95 ;
		RECT	0 29.25 0.32 29.61 ;
		RECT	0 30.31 0.32 31.95 ;
		RECT	0 32.555 0.32 32.77 ;
		RECT	0 33.07 0.32 33.175 ;
		RECT	0 33.475 0.32 35.285 ;
		RECT	0 35.585 0.32 35.8 ;
		RECT	0 36.1 0.32 36.205 ;
		RECT	0 36.505 0.32 36.94 ;
		RECT	0 37.24 0.32 37.345 ;
		RECT	0 37.645 0.32 37.86 ;
		RECT	0 38.16 0.32 38.345 ;
		RECT	0 38.645 0.32 38.83 ;
		RECT	0 39.13 0.32 39.235 ;
		RECT	0 39.535 0.32 39.63 ;
		RECT	0 39.93 0.32 40 ;
		RECT	0 40.3 0.32 40.375 ;
		RECT	0 40.675 0.32 40.86 ;
		RECT	0 41.77 0.32 41.86 ;
		RECT	0 42.16 0.32 42.265 ;
		RECT	0 42.565 0.32 43.005 ;
		RECT	0 43.705 0.32 43.89 ;
		RECT	0 44.705 0.32 44.89 ;
		RECT	0 45.19 0.32 45.295 ;
		RECT	0 45.595 0.32 47.4 ;
		RECT	0 48.1 0.32 48.57 ;
		RECT	0 48.87 0.32 50.235 ;
		RECT	0 50.535 0.32 53.16 ;
		RECT	0 53.46 0.32 53.565 ;
		RECT	0 53.865 0.32 54.05 ;
		RECT	0 54.86 0.32 55.05 ;
		RECT	0 55.35 0.32 55.425 ;
		RECT	0 55.725 0.32 55.805 ;
		RECT	0 56.105 0.32 56.19 ;
		RECT	0 56.49 0.32 56.595 ;
		RECT	0 57.38 0.32 57.595 ;
		RECT	0 57.895 0.32 58.08 ;
		RECT	0 58.38 0.32 58.485 ;
		RECT	0 58.785 0.32 59.25 ;
		RECT	0 59.55 0.32 59.625 ;
		RECT	0 59.925 0.32 60.08 ;
		RECT	0 60.925 0.32 61.11 ;
		RECT	0 61.41 0.32 61.485 ;
		RECT	0 62.125 0.32 62.25 ;
		RECT	0 62.76 0.32 63.14 ;
		RECT	0 63.44 0.32 65.28 ;
		RECT	0 65.58 0.32 65.685 ;
		RECT	0 65.985 0.32 66.17 ;
		RECT	0 66.725 0.32 67.2 ;
		RECT	0 67.5 0.32 69.81 ;
		RECT	0 70.11 0.32 70.205 ;
		RECT	0 70.505 0.32 70.75 ;
		RECT	0 71.05 0.32 72.365 ;
		RECT	0 72.925 0.32 73.355 ;
		RECT	0 73.655 0.32 75.245 ;
		RECT	0 75.805 0.32 76.235 ;
		RECT	0 76.535 0.32 78.125 ;
		RECT	0 78.685 0.32 79.115 ;
		RECT	0 79.415 0.32 81.005 ;
		RECT	0 81.565 0.32 81.995 ;
		RECT	0 82.295 0.32 83.885 ;
		RECT	0 84.445 0.32 84.875 ;
		RECT	0 85.175 0.32 86.765 ;
		RECT	0 87.325 0.32 87.755 ;
		RECT	0 88.055 0.32 89.645 ;
		RECT	0 90.205 0.32 90.635 ;
		RECT	0 90.935 0.32 92.525 ;
		RECT	0 93.085 0.32 93.515 ;
		RECT	0 93.815 0.32 95.405 ;
		RECT	0 95.965 0.32 96.395 ;
		RECT	0 96.695 0.32 98.285 ;
		RECT	0 98.845 0.32 99.275 ;
		RECT	0 99.575 0.32 100.38 ;
		RECT	51.085 0 51.405 100.94 ;
		RECT	0.32 0 51.085 0.35 ;
		RECT	0.32 100.59 51.085 100.94 ;
		LAYER	M3 DESIGNRULEWIDTH 0.165 ;
		RECT	0.32 0.35 51.085 100.59 ;
		RECT	0 0.56 0.32 1.365 ;
		RECT	0 1.665 0.32 2.095 ;
		RECT	0 2.655 0.32 4.245 ;
		RECT	0 4.545 0.32 4.975 ;
		RECT	0 5.535 0.32 7.125 ;
		RECT	0 7.425 0.32 7.855 ;
		RECT	0 8.415 0.32 10.005 ;
		RECT	0 10.305 0.32 10.735 ;
		RECT	0 11.295 0.32 12.885 ;
		RECT	0 13.185 0.32 13.615 ;
		RECT	0 14.175 0.32 15.765 ;
		RECT	0 16.065 0.32 16.495 ;
		RECT	0 17.055 0.32 18.645 ;
		RECT	0 18.945 0.32 19.375 ;
		RECT	0 19.935 0.32 21.525 ;
		RECT	0 21.825 0.32 22.255 ;
		RECT	0 22.815 0.32 24.405 ;
		RECT	0 24.705 0.32 25.135 ;
		RECT	0 25.695 0.32 28.6 ;
		RECT	0 28.9 0.32 28.95 ;
		RECT	0 29.25 0.32 29.61 ;
		RECT	0 30.31 0.32 31.95 ;
		RECT	0 32.555 0.32 32.77 ;
		RECT	0 33.07 0.32 33.175 ;
		RECT	0 33.475 0.32 35.285 ;
		RECT	0 35.585 0.32 35.8 ;
		RECT	0 36.1 0.32 36.205 ;
		RECT	0 36.505 0.32 36.94 ;
		RECT	0 37.24 0.32 37.345 ;
		RECT	0 37.645 0.32 37.86 ;
		RECT	0 38.16 0.32 38.345 ;
		RECT	0 38.645 0.32 38.83 ;
		RECT	0 39.13 0.32 39.235 ;
		RECT	0 39.535 0.32 39.63 ;
		RECT	0 39.93 0.32 40 ;
		RECT	0 40.3 0.32 40.375 ;
		RECT	0 40.675 0.32 40.86 ;
		RECT	0 41.77 0.32 41.86 ;
		RECT	0 42.16 0.32 42.265 ;
		RECT	0 42.565 0.32 43.005 ;
		RECT	0 43.705 0.32 43.89 ;
		RECT	0 44.705 0.32 44.89 ;
		RECT	0 45.19 0.32 45.295 ;
		RECT	0 45.595 0.32 47.4 ;
		RECT	0 48.1 0.32 48.57 ;
		RECT	0 48.87 0.32 50.235 ;
		RECT	0 50.535 0.32 53.16 ;
		RECT	0 53.46 0.32 53.565 ;
		RECT	0 53.865 0.32 54.05 ;
		RECT	0 54.86 0.32 55.05 ;
		RECT	0 55.35 0.32 55.425 ;
		RECT	0 55.725 0.32 55.805 ;
		RECT	0 56.105 0.32 56.19 ;
		RECT	0 56.49 0.32 56.595 ;
		RECT	0 57.38 0.32 57.595 ;
		RECT	0 57.895 0.32 58.08 ;
		RECT	0 58.38 0.32 58.485 ;
		RECT	0 58.785 0.32 59.25 ;
		RECT	0 59.55 0.32 59.625 ;
		RECT	0 59.925 0.32 60.08 ;
		RECT	0 60.925 0.32 61.11 ;
		RECT	0 61.41 0.32 61.485 ;
		RECT	0 62.125 0.32 62.25 ;
		RECT	0 62.76 0.32 63.14 ;
		RECT	0 63.44 0.32 65.28 ;
		RECT	0 65.58 0.32 65.685 ;
		RECT	0 65.985 0.32 66.17 ;
		RECT	0 66.725 0.32 67.2 ;
		RECT	0 67.5 0.32 69.81 ;
		RECT	0 70.11 0.32 70.205 ;
		RECT	0 70.505 0.32 70.75 ;
		RECT	0 71.05 0.32 72.365 ;
		RECT	0 72.925 0.32 73.355 ;
		RECT	0 73.655 0.32 75.245 ;
		RECT	0 75.805 0.32 76.235 ;
		RECT	0 76.535 0.32 78.125 ;
		RECT	0 78.685 0.32 79.115 ;
		RECT	0 79.415 0.32 81.005 ;
		RECT	0 81.565 0.32 81.995 ;
		RECT	0 82.295 0.32 83.885 ;
		RECT	0 84.445 0.32 84.875 ;
		RECT	0 85.175 0.32 86.765 ;
		RECT	0 87.325 0.32 87.755 ;
		RECT	0 88.055 0.32 89.645 ;
		RECT	0 90.205 0.32 90.635 ;
		RECT	0 90.935 0.32 92.525 ;
		RECT	0 93.085 0.32 93.515 ;
		RECT	0 93.815 0.32 95.405 ;
		RECT	0 95.965 0.32 96.395 ;
		RECT	0 96.695 0.32 98.285 ;
		RECT	0 98.845 0.32 99.275 ;
		RECT	0 99.575 0.32 100.38 ;
		RECT	51.085 0 51.405 100.94 ;
		RECT	0.32 0 51.085 0.35 ;
		RECT	0.32 100.59 51.085 100.94 ;
		LAYER	M4 DESIGNRULEWIDTH 0.165 ;
		RECT	0.57 26.775 14.49 27.945 ;
		RECT	14.185 27.945 14.49 28.175 ;
		RECT	0.57 28.005 14.125 28.155 ;
		RECT	0.57 28.905 14.49 29.015 ;
		RECT	0.57 29.15 14.49 29.34 ;
		RECT	0.57 29.825 14.49 29.925 ;
		RECT	0.57 30.315 11.56 30.415 ;
		RECT	0.57 30.805 14.49 30.905 ;
		RECT	11.255 30.905 14.49 30.91 ;
		RECT	11.255 30.91 12.345 31.255 ;
		RECT	0.57 31.005 11.155 31.215 ;
		RECT	12.445 31.01 14.49 31.2 ;
		RECT	11.255 31.255 11.56 31.315 ;
		RECT	0.57 31.315 11.56 31.385 ;
		RECT	0.57 31.485 14.49 31.675 ;
		RECT	0.57 31.775 14.49 31.93 ;
		RECT	0.57 32.32 14.49 32.385 ;
		RECT	0.57 32.775 14.49 32.88 ;
		RECT	0.57 33.27 14.49 33.37 ;
		RECT	0.57 33.76 14.15 33.86 ;
		RECT	0.57 34.25 14.49 34.355 ;
		RECT	0.57 34.745 14.49 34.845 ;
		RECT	0.57 35.235 14.49 35.34 ;
		RECT	0.57 35.44 14.49 35.63 ;
		RECT	0.57 35.73 14.49 35.83 ;
		RECT	0.57 36.22 14.49 36.325 ;
		RECT	0.57 36.715 14.49 36.815 ;
		RECT	0.57 37.205 14.49 37.305 ;
		RECT	0.57 37.695 14.49 37.8 ;
		RECT	0.57 38.19 14.49 38.29 ;
		RECT	0.57 38.68 14.49 38.78 ;
		RECT	0.57 39.17 14.49 39.275 ;
		RECT	0.57 39.375 14.49 39.565 ;
		RECT	0.57 39.665 14.49 39.765 ;
		RECT	0.57 40.155 14.49 40.26 ;
		RECT	0.57 40.65 14.49 40.75 ;
		RECT	8.61 41.14 14.49 41.23 ;
		RECT	0.57 41.155 8.56 41.225 ;
		RECT	0.57 41.64 14.49 41.735 ;
		RECT	0.57 42.125 14.49 42.225 ;
		RECT	0.57 42.615 14.49 42.72 ;
		RECT	9.515 43.11 14.49 43.2 ;
		RECT	9.295 43.115 9.465 43.125 ;
		RECT	0.57 43.125 9.465 43.195 ;
		RECT	9.295 43.195 9.465 43.205 ;
		RECT	0.57 43.3 14.49 43.51 ;
		RECT	0.57 43.61 14.49 43.705 ;
		RECT	0.57 44.095 14.49 44.2 ;
		RECT	0.57 44.59 14.49 44.685 ;
		RECT	0.57 45.075 14.49 45.18 ;
		RECT	0.57 45.57 14.49 45.655 ;
		RECT	0.57 46.045 14.49 46.28 ;
		RECT	0.57 46.28 13.465 46.395 ;
		RECT	13.565 46.38 14.49 46.57 ;
		RECT	11.215 46.395 13.465 46.655 ;
		RECT	0.57 46.455 11.155 46.605 ;
		RECT	0.57 47.045 13.8 47.145 ;
		RECT	0.57 47.245 14.49 47.435 ;
		RECT	0.57 47.535 13.8 47.64 ;
		RECT	0.57 48.03 14.49 48.13 ;
		RECT	0.57 48.52 14.49 48.62 ;
		RECT	0.57 49.01 7.02 49.115 ;
		RECT	13.595 49.01 14.49 49.115 ;
		RECT	0.57 49.505 14.49 49.605 ;
		RECT	0.57 49.995 14.49 50.1 ;
		RECT	0.57 50.49 13.8 50.59 ;
		RECT	0.57 50.69 14.49 50.88 ;
		RECT	0.57 50.98 13.8 51.08 ;
		RECT	11.215 51.47 13.5 51.73 ;
		RECT	13.6 51.495 14.49 51.685 ;
		RECT	0.57 51.52 11.155 51.67 ;
		RECT	0.57 51.73 13.5 51.785 ;
		RECT	0.57 51.785 14.49 52.08 ;
		RECT	0.57 52.47 14.49 52.555 ;
		RECT	0.57 52.945 14.49 53.05 ;
		RECT	0.57 53.44 14.49 53.545 ;
		RECT	0.57 53.935 14.49 54.025 ;
		RECT	7.785 54.435 14.49 54.515 ;
		RECT	0.57 54.44 7.735 54.51 ;
		RECT	0.57 54.615 14.49 54.825 ;
		RECT	0.57 54.925 14.49 55.02 ;
		RECT	0.57 55.41 14.49 55.51 ;
		RECT	0.57 55.9 14.49 56.005 ;
		RECT	0.57 56.395 14.49 56.485 ;
		RECT	8.06 56.895 14.49 56.985 ;
		RECT	0.57 56.9 8.01 56.97 ;
		RECT	0.57 57.375 14.49 57.48 ;
		RECT	0.57 57.87 14.49 57.97 ;
		RECT	0.57 58.36 14.49 58.465 ;
		RECT	0.57 58.565 14.49 58.755 ;
		RECT	0.57 58.855 14.49 58.955 ;
		RECT	0.57 59.345 14.49 59.445 ;
		RECT	0.57 59.835 14.49 59.94 ;
		RECT	0.57 60.33 14.49 60.43 ;
		RECT	0.57 60.82 14.49 60.925 ;
		RECT	0.57 61.315 14.49 61.415 ;
		RECT	0.57 61.805 14.49 61.905 ;
		RECT	0.57 62.295 14.15 62.39 ;
		RECT	0.57 62.49 14.49 62.7 ;
		RECT	2.785 62.8 14.49 62.89 ;
		RECT	0.57 63.28 14.49 63.375 ;
		RECT	0.57 63.79 14.49 63.86 ;
		RECT	0.57 64.28 14.49 64.35 ;
		RECT	0.57 64.765 14.49 64.825 ;
		RECT	0.57 65.215 14.49 65.35 ;
		RECT	0.57 65.74 14.49 65.81 ;
		RECT	0.57 66.2 14.49 66.35 ;
		RECT	0.57 66.45 14.49 66.64 ;
		RECT	0.57 66.74 12.555 66.815 ;
		RECT	11.255 66.815 12.555 66.825 ;
		RECT	11.255 66.825 12.27 67.215 ;
		RECT	0.57 66.915 11.155 67.125 ;
		RECT	12.37 66.925 14.49 67.115 ;
		RECT	11.255 67.215 14.49 67.225 ;
		RECT	0.57 67.225 14.49 67.32 ;
		RECT	0.57 67.71 12.555 67.81 ;
		RECT	0.57 68.2 14.49 68.305 ;
		RECT	0.57 68.705 14.49 68.915 ;
		RECT	0.57 69.045 14.49 69.155 ;
		RECT	14.21 69.885 14.49 70.115 ;
		RECT	0.57 69.905 14.15 70.055 ;
		RECT	0.57 70.115 14.49 71.285 ;
		RECT	0.21 28.005 0.57 28.155 ;
		RECT	0.215 29.15 0.57 29.34 ;
		RECT	0.22 31.005 0.57 31.215 ;
		RECT	0.22 31.485 0.57 31.675 ;
		RECT	0.22 35.44 0.57 35.63 ;
		RECT	0.23 39.375 0.57 39.565 ;
		RECT	0.14 41.155 0.57 41.225 ;
		RECT	0.15 43.125 0.57 43.195 ;
		RECT	0.215 43.3 0.57 43.51 ;
		RECT	0.21 46.455 0.57 46.605 ;
		RECT	0.225 47.245 0.57 47.435 ;
		RECT	0.325 50.69 0.61 50.88 ;
		RECT	0.21 51.52 0.57 51.67 ;
		RECT	0.15 54.44 0.57 54.51 ;
		RECT	0.235 54.615 0.57 54.825 ;
		RECT	0.14 56.9 0.57 56.97 ;
		RECT	0.24 58.565 0.57 58.755 ;
		RECT	0.225 62.49 0.57 62.7 ;
		RECT	0.14 62.805 0.57 62.875 ;
		RECT	0.235 66.45 0.57 66.64 ;
		RECT	0.225 66.915 0.57 67.125 ;
		RECT	0.24 68.705 0.57 68.915 ;
		RECT	0.22 69.905 0.57 70.055 ;
		RECT	5.7 23.225 13.945 23.375 ;
		RECT	5.7 20.345 13.945 20.495 ;
		RECT	5.7 17.465 13.945 17.615 ;
		RECT	5.7 14.585 13.945 14.735 ;
		RECT	5.7 11.705 13.945 11.855 ;
		RECT	5.7 8.825 13.945 8.975 ;
		RECT	5.7 5.945 13.945 6.095 ;
		RECT	5.7 3.065 13.945 3.215 ;
		RECT	5.7 26.105 13.945 26.255 ;
		RECT	0.57 23.225 1.11 23.375 ;
		RECT	0.57 20.345 1.11 20.495 ;
		RECT	0.57 17.465 1.11 17.615 ;
		RECT	0.57 14.585 1.11 14.735 ;
		RECT	0.57 11.705 1.11 11.855 ;
		RECT	0.57 8.825 1.11 8.975 ;
		RECT	0.57 5.945 1.11 6.095 ;
		RECT	0.57 3.065 1.11 3.215 ;
		RECT	0.57 26.105 1.11 26.255 ;
		RECT	1.005 23.225 5.7 23.375 ;
		RECT	1.005 20.345 5.7 20.495 ;
		RECT	1.005 17.465 5.7 17.615 ;
		RECT	1.005 14.585 5.7 14.735 ;
		RECT	1.005 11.705 5.7 11.855 ;
		RECT	1.005 8.825 5.7 8.975 ;
		RECT	1.005 5.945 5.7 6.095 ;
		RECT	1.005 3.065 5.7 3.215 ;
		RECT	1.005 26.105 5.7 26.255 ;
		RECT	0.255 26.105 0.57 26.255 ;
		RECT	0.255 23.225 0.57 23.375 ;
		RECT	0.255 20.345 0.57 20.495 ;
		RECT	0.255 17.465 0.57 17.615 ;
		RECT	0.255 14.585 0.57 14.735 ;
		RECT	0.255 11.705 0.57 11.855 ;
		RECT	0.255 8.825 0.57 8.975 ;
		RECT	0.255 5.945 0.57 6.095 ;
		RECT	0.255 3.065 0.57 3.215 ;
		RECT	5.7 74.685 13.945 74.835 ;
		RECT	5.7 77.565 13.945 77.715 ;
		RECT	5.7 80.445 13.945 80.595 ;
		RECT	5.7 83.325 13.945 83.475 ;
		RECT	5.7 86.205 13.945 86.355 ;
		RECT	5.7 89.085 13.945 89.235 ;
		RECT	5.7 91.965 13.945 92.115 ;
		RECT	5.7 94.845 13.945 94.995 ;
		RECT	5.7 97.725 13.945 97.875 ;
		RECT	5.7 71.805 13.945 71.955 ;
		RECT	0.57 74.685 1.11 74.835 ;
		RECT	0.57 77.565 1.11 77.715 ;
		RECT	0.57 80.445 1.11 80.595 ;
		RECT	0.57 83.325 1.11 83.475 ;
		RECT	0.57 86.205 1.11 86.355 ;
		RECT	0.57 89.085 1.11 89.235 ;
		RECT	0.57 91.965 1.11 92.115 ;
		RECT	0.57 94.845 1.11 94.995 ;
		RECT	0.57 97.725 1.11 97.875 ;
		RECT	0.57 71.805 1.11 71.955 ;
		RECT	1.005 74.685 5.7 74.835 ;
		RECT	1.005 77.565 5.7 77.715 ;
		RECT	1.005 80.445 5.7 80.595 ;
		RECT	1.005 83.325 5.7 83.475 ;
		RECT	1.005 86.205 5.7 86.355 ;
		RECT	1.005 89.085 5.7 89.235 ;
		RECT	1.005 91.965 5.7 92.115 ;
		RECT	1.005 94.845 5.7 94.995 ;
		RECT	1.005 97.725 5.7 97.875 ;
		RECT	1.005 71.805 5.7 71.955 ;
		RECT	0.255 71.805 0.57 71.955 ;
		RECT	0.255 74.685 0.57 74.835 ;
		RECT	0.255 77.565 0.57 77.715 ;
		RECT	0.255 80.445 0.57 80.595 ;
		RECT	0.255 83.325 0.57 83.475 ;
		RECT	0.255 86.205 0.57 86.355 ;
		RECT	0.255 89.085 0.57 89.235 ;
		RECT	0.255 91.965 0.57 92.115 ;
		RECT	0.255 94.845 0.57 94.995 ;
		RECT	0.255 97.725 0.57 97.875 ;
		RECT	15.63 28.905 16.17 29.015 ;
		RECT	15.63 26.775 16.17 28.175 ;
		RECT	16.17 28.905 16.71 29.015 ;
		RECT	16.17 26.775 16.71 28.175 ;
		RECT	16.71 28.905 17.25 29.015 ;
		RECT	16.71 26.775 17.25 28.175 ;
		RECT	15.09 28.905 15.63 29.015 ;
		RECT	15.09 26.775 15.63 28.175 ;
		RECT	14.49 28.905 15.09 29.015 ;
		RECT	14.49 26.775 15.09 28.175 ;
		RECT	19.41 28.905 19.95 29.015 ;
		RECT	19.41 26.775 19.95 28.175 ;
		RECT	19.95 28.905 20.49 29.015 ;
		RECT	19.95 26.775 20.49 28.175 ;
		RECT	20.49 28.905 21.03 29.015 ;
		RECT	20.49 26.775 21.03 28.175 ;
		RECT	21.03 28.905 21.57 29.015 ;
		RECT	21.03 26.775 21.57 28.175 ;
		RECT	21.57 28.905 22.11 29.015 ;
		RECT	21.57 26.775 22.11 28.175 ;
		RECT	22.11 28.905 22.65 29.015 ;
		RECT	22.11 26.775 22.65 28.175 ;
		RECT	22.65 28.905 23.19 29.015 ;
		RECT	22.65 26.775 23.19 28.175 ;
		RECT	23.19 28.905 23.73 29.015 ;
		RECT	23.19 26.775 23.73 28.175 ;
		RECT	23.73 28.905 24.27 29.015 ;
		RECT	23.73 26.775 24.27 28.175 ;
		RECT	24.27 28.905 24.81 29.015 ;
		RECT	24.27 26.775 24.81 28.175 ;
		RECT	24.81 28.905 25.35 29.015 ;
		RECT	24.81 26.775 25.35 28.175 ;
		RECT	25.35 28.905 25.89 29.015 ;
		RECT	25.35 26.775 25.89 28.175 ;
		RECT	25.89 28.905 26.43 29.015 ;
		RECT	25.89 26.775 26.43 28.175 ;
		RECT	26.43 28.905 26.97 29.015 ;
		RECT	26.43 26.775 26.97 28.175 ;
		RECT	26.97 28.905 27.51 29.015 ;
		RECT	26.97 26.775 27.51 28.175 ;
		RECT	27.51 28.905 28.05 29.015 ;
		RECT	27.51 26.775 28.05 28.175 ;
		RECT	28.05 28.905 28.59 29.015 ;
		RECT	28.05 26.775 28.59 28.175 ;
		RECT	28.59 28.905 29.13 29.015 ;
		RECT	28.59 26.775 29.13 28.175 ;
		RECT	29.13 28.905 29.67 29.015 ;
		RECT	29.13 26.775 29.67 28.175 ;
		RECT	29.67 28.905 30.21 29.015 ;
		RECT	29.67 26.775 30.21 28.175 ;
		RECT	30.21 28.905 30.75 29.015 ;
		RECT	30.21 26.775 30.75 28.175 ;
		RECT	30.75 28.905 31.29 29.015 ;
		RECT	30.75 26.775 31.29 28.175 ;
		RECT	31.29 28.905 31.83 29.015 ;
		RECT	31.29 26.775 31.83 28.175 ;
		RECT	31.83 28.905 32.37 29.015 ;
		RECT	31.83 26.775 32.37 28.175 ;
		RECT	32.37 28.905 32.91 29.015 ;
		RECT	32.37 26.775 32.91 28.175 ;
		RECT	32.91 28.905 33.45 29.015 ;
		RECT	32.91 26.775 33.45 28.175 ;
		RECT	33.45 28.905 33.99 29.015 ;
		RECT	33.45 26.775 33.99 28.175 ;
		RECT	33.99 28.905 34.53 29.015 ;
		RECT	33.99 26.775 34.53 28.175 ;
		RECT	34.53 28.905 35.07 29.015 ;
		RECT	34.53 26.775 35.07 28.175 ;
		RECT	35.07 28.905 35.61 29.015 ;
		RECT	35.07 26.775 35.61 28.175 ;
		RECT	35.61 28.905 36.15 29.015 ;
		RECT	35.61 26.775 36.15 28.175 ;
		RECT	36.15 28.905 36.69 29.015 ;
		RECT	36.15 26.775 36.69 28.175 ;
		RECT	36.69 28.905 37.23 29.015 ;
		RECT	36.69 26.775 37.23 28.175 ;
		RECT	37.23 28.905 37.77 29.015 ;
		RECT	37.23 26.775 37.77 28.175 ;
		RECT	37.77 28.905 38.31 29.015 ;
		RECT	37.77 26.775 38.31 28.175 ;
		RECT	38.31 28.905 38.85 29.015 ;
		RECT	38.31 26.775 38.85 28.175 ;
		RECT	38.85 28.905 39.39 29.015 ;
		RECT	38.85 26.775 39.39 28.175 ;
		RECT	39.39 28.905 39.93 29.015 ;
		RECT	39.39 26.775 39.93 28.175 ;
		RECT	39.93 28.905 40.47 29.015 ;
		RECT	39.93 26.775 40.47 28.175 ;
		RECT	40.47 28.905 41.01 29.015 ;
		RECT	40.47 26.775 41.01 28.175 ;
		RECT	41.01 28.905 41.55 29.015 ;
		RECT	41.01 26.775 41.55 28.175 ;
		RECT	41.55 28.905 42.09 29.015 ;
		RECT	41.55 26.775 42.09 28.175 ;
		RECT	42.09 28.905 42.63 29.015 ;
		RECT	42.09 26.775 42.63 28.175 ;
		RECT	42.63 28.905 43.17 29.015 ;
		RECT	42.63 26.775 43.17 28.175 ;
		RECT	43.17 28.905 43.71 29.015 ;
		RECT	43.17 26.775 43.71 28.175 ;
		RECT	43.71 28.905 44.25 29.015 ;
		RECT	43.71 26.775 44.25 28.175 ;
		RECT	44.25 28.905 44.79 29.015 ;
		RECT	44.25 26.775 44.79 28.175 ;
		RECT	44.79 28.905 45.33 29.015 ;
		RECT	44.79 26.775 45.33 28.175 ;
		RECT	45.33 28.905 45.87 29.015 ;
		RECT	45.33 26.775 45.87 28.175 ;
		RECT	45.87 28.905 46.41 29.015 ;
		RECT	45.87 26.775 46.41 28.175 ;
		RECT	17.25 28.905 17.79 29.015 ;
		RECT	17.25 26.775 17.79 28.175 ;
		RECT	46.41 28.905 46.95 29.015 ;
		RECT	46.41 26.775 46.95 28.175 ;
		RECT	46.95 28.905 47.49 29.015 ;
		RECT	46.95 26.775 47.49 28.175 ;
		RECT	47.49 28.905 48.03 29.015 ;
		RECT	47.49 26.775 48.03 28.175 ;
		RECT	48.03 28.905 48.57 29.015 ;
		RECT	48.03 26.775 48.57 28.175 ;
		RECT	48.57 28.905 49.11 29.015 ;
		RECT	48.57 26.775 49.11 28.175 ;
		RECT	17.79 28.905 18.33 29.015 ;
		RECT	17.79 26.775 18.33 28.175 ;
		RECT	18.33 28.905 18.87 29.015 ;
		RECT	18.33 26.775 18.87 28.175 ;
		RECT	18.87 28.905 19.41 29.015 ;
		RECT	18.87 26.775 19.41 28.175 ;
		RECT	49.65 28.905 50.25 29.015 ;
		RECT	49.65 26.775 50.25 28.175 ;
		RECT	49.11 28.905 49.65 29.015 ;
		RECT	49.11 26.775 49.65 28.175 ;
		RECT	15.09 69.045 15.63 69.155 ;
		RECT	15.09 69.885 15.63 71.285 ;
		RECT	14.49 69.045 15.09 69.155 ;
		RECT	14.49 69.885 15.09 71.285 ;
		RECT	19.41 69.045 19.95 69.155 ;
		RECT	19.41 69.885 19.95 71.285 ;
		RECT	19.95 69.045 20.49 69.155 ;
		RECT	19.95 69.885 20.49 71.285 ;
		RECT	20.49 69.045 21.03 69.155 ;
		RECT	20.49 69.885 21.03 71.285 ;
		RECT	21.03 69.045 21.57 69.155 ;
		RECT	21.03 69.885 21.57 71.285 ;
		RECT	21.57 69.045 22.11 69.155 ;
		RECT	21.57 69.885 22.11 71.285 ;
		RECT	22.11 69.045 22.65 69.155 ;
		RECT	22.11 69.885 22.65 71.285 ;
		RECT	22.65 69.045 23.19 69.155 ;
		RECT	22.65 69.885 23.19 71.285 ;
		RECT	23.19 69.045 23.73 69.155 ;
		RECT	23.19 69.885 23.73 71.285 ;
		RECT	23.73 69.045 24.27 69.155 ;
		RECT	23.73 69.885 24.27 71.285 ;
		RECT	24.27 69.045 24.81 69.155 ;
		RECT	24.27 69.885 24.81 71.285 ;
		RECT	24.81 69.045 25.35 69.155 ;
		RECT	24.81 69.885 25.35 71.285 ;
		RECT	25.35 69.045 25.89 69.155 ;
		RECT	25.35 69.885 25.89 71.285 ;
		RECT	25.89 69.045 26.43 69.155 ;
		RECT	25.89 69.885 26.43 71.285 ;
		RECT	26.43 69.045 26.97 69.155 ;
		RECT	26.43 69.885 26.97 71.285 ;
		RECT	26.97 69.045 27.51 69.155 ;
		RECT	26.97 69.885 27.51 71.285 ;
		RECT	27.51 69.045 28.05 69.155 ;
		RECT	27.51 69.885 28.05 71.285 ;
		RECT	28.05 69.045 28.59 69.155 ;
		RECT	28.05 69.885 28.59 71.285 ;
		RECT	28.59 69.045 29.13 69.155 ;
		RECT	28.59 69.885 29.13 71.285 ;
		RECT	29.13 69.045 29.67 69.155 ;
		RECT	29.13 69.885 29.67 71.285 ;
		RECT	29.67 69.045 30.21 69.155 ;
		RECT	29.67 69.885 30.21 71.285 ;
		RECT	15.63 69.045 16.17 69.155 ;
		RECT	15.63 69.885 16.17 71.285 ;
		RECT	30.21 69.045 30.75 69.155 ;
		RECT	30.21 69.885 30.75 71.285 ;
		RECT	30.75 69.045 31.29 69.155 ;
		RECT	30.75 69.885 31.29 71.285 ;
		RECT	31.29 69.045 31.83 69.155 ;
		RECT	31.29 69.885 31.83 71.285 ;
		RECT	31.83 69.045 32.37 69.155 ;
		RECT	31.83 69.885 32.37 71.285 ;
		RECT	32.37 69.045 32.91 69.155 ;
		RECT	32.37 69.885 32.91 71.285 ;
		RECT	32.91 69.045 33.45 69.155 ;
		RECT	32.91 69.885 33.45 71.285 ;
		RECT	33.45 69.045 33.99 69.155 ;
		RECT	33.45 69.885 33.99 71.285 ;
		RECT	33.99 69.045 34.53 69.155 ;
		RECT	33.99 69.885 34.53 71.285 ;
		RECT	34.53 69.045 35.07 69.155 ;
		RECT	34.53 69.885 35.07 71.285 ;
		RECT	35.07 69.045 35.61 69.155 ;
		RECT	35.07 69.885 35.61 71.285 ;
		RECT	16.17 69.045 16.71 69.155 ;
		RECT	16.17 69.885 16.71 71.285 ;
		RECT	35.61 69.045 36.15 69.155 ;
		RECT	35.61 69.885 36.15 71.285 ;
		RECT	36.15 69.045 36.69 69.155 ;
		RECT	36.15 69.885 36.69 71.285 ;
		RECT	36.69 69.045 37.23 69.155 ;
		RECT	36.69 69.885 37.23 71.285 ;
		RECT	37.23 69.045 37.77 69.155 ;
		RECT	37.23 69.885 37.77 71.285 ;
		RECT	37.77 69.045 38.31 69.155 ;
		RECT	37.77 69.885 38.31 71.285 ;
		RECT	38.31 69.045 38.85 69.155 ;
		RECT	38.31 69.885 38.85 71.285 ;
		RECT	38.85 69.045 39.39 69.155 ;
		RECT	38.85 69.885 39.39 71.285 ;
		RECT	39.39 69.045 39.93 69.155 ;
		RECT	39.39 69.885 39.93 71.285 ;
		RECT	39.93 69.045 40.47 69.155 ;
		RECT	39.93 69.885 40.47 71.285 ;
		RECT	40.47 69.045 41.01 69.155 ;
		RECT	40.47 69.885 41.01 71.285 ;
		RECT	16.71 69.045 17.25 69.155 ;
		RECT	16.71 69.885 17.25 71.285 ;
		RECT	41.01 69.045 41.55 69.155 ;
		RECT	41.01 69.885 41.55 71.285 ;
		RECT	41.55 69.045 42.09 69.155 ;
		RECT	41.55 69.885 42.09 71.285 ;
		RECT	42.09 69.045 42.63 69.155 ;
		RECT	42.09 69.885 42.63 71.285 ;
		RECT	42.63 69.045 43.17 69.155 ;
		RECT	42.63 69.885 43.17 71.285 ;
		RECT	43.17 69.045 43.71 69.155 ;
		RECT	43.17 69.885 43.71 71.285 ;
		RECT	43.71 69.045 44.25 69.155 ;
		RECT	43.71 69.885 44.25 71.285 ;
		RECT	44.25 69.045 44.79 69.155 ;
		RECT	44.25 69.885 44.79 71.285 ;
		RECT	44.79 69.045 45.33 69.155 ;
		RECT	44.79 69.885 45.33 71.285 ;
		RECT	45.33 69.045 45.87 69.155 ;
		RECT	45.33 69.885 45.87 71.285 ;
		RECT	45.87 69.045 46.41 69.155 ;
		RECT	45.87 69.885 46.41 71.285 ;
		RECT	17.25 69.045 17.79 69.155 ;
		RECT	17.25 69.885 17.79 71.285 ;
		RECT	46.41 69.045 46.95 69.155 ;
		RECT	46.41 69.885 46.95 71.285 ;
		RECT	46.95 69.045 47.49 69.155 ;
		RECT	46.95 69.885 47.49 71.285 ;
		RECT	47.49 69.045 48.03 69.155 ;
		RECT	47.49 69.885 48.03 71.285 ;
		RECT	48.03 69.045 48.57 69.155 ;
		RECT	48.03 69.885 48.57 71.285 ;
		RECT	48.57 69.045 49.11 69.155 ;
		RECT	48.57 69.885 49.11 71.285 ;
		RECT	17.79 69.045 18.33 69.155 ;
		RECT	17.79 69.885 18.33 71.285 ;
		RECT	18.33 69.045 18.87 69.155 ;
		RECT	18.33 69.885 18.87 71.285 ;
		RECT	18.87 69.045 19.41 69.155 ;
		RECT	18.87 69.885 19.41 71.285 ;
		RECT	49.65 69.045 50.25 69.155 ;
		RECT	49.65 69.885 50.25 71.285 ;
		RECT	49.11 69.045 49.65 69.155 ;
		RECT	49.11 69.885 49.65 71.285 ;
		RECT	50.25 26.775 51.405 28.175 ;
		RECT	50.25 28.905 51.405 29.015 ;
		RECT	51.21 29.015 51.405 29.435 ;
		RECT	50.25 29.15 51.11 29.34 ;
		RECT	50.25 29.825 51.405 29.925 ;
		RECT	50.25 30.805 51.405 30.91 ;
		RECT	51.21 30.91 51.405 31.255 ;
		RECT	50.25 31.01 51.11 31.2 ;
		RECT	51.21 31.435 51.405 31.775 ;
		RECT	50.25 31.485 51.11 31.675 ;
		RECT	51.16 31.775 51.405 31.93 ;
		RECT	50.25 31.78 51.1 31.93 ;
		RECT	50.25 32.32 51.405 32.385 ;
		RECT	50.25 32.775 51.405 32.88 ;
		RECT	50.25 33.27 51.405 33.37 ;
		RECT	50.65 33.76 51.405 33.86 ;
		RECT	50.25 34.25 51.405 34.355 ;
		RECT	51.03 34.355 51.405 34.745 ;
		RECT	50.25 34.745 51.405 34.845 ;
		RECT	50.25 35.235 51.405 35.34 ;
		RECT	51.21 35.34 51.405 35.73 ;
		RECT	50.25 35.44 51.11 35.63 ;
		RECT	50.25 35.73 51.405 35.83 ;
		RECT	50.25 36.22 51.405 36.325 ;
		RECT	50.25 36.715 51.405 36.815 ;
		RECT	50.25 37.205 51.405 37.305 ;
		RECT	50.25 37.695 51.405 37.8 ;
		RECT	50.25 38.19 51.405 38.29 ;
		RECT	50.25 38.68 51.405 38.78 ;
		RECT	50.25 39.17 51.405 39.275 ;
		RECT	51.21 39.275 51.405 39.665 ;
		RECT	50.25 39.375 51.11 39.565 ;
		RECT	50.25 39.665 51.405 39.765 ;
		RECT	50.25 40.155 51.405 40.26 ;
		RECT	50.25 40.65 51.405 40.75 ;
		RECT	50.25 41.14 51.405 41.23 ;
		RECT	50.25 41.64 51.405 41.735 ;
		RECT	50.25 42.125 51.405 42.225 ;
		RECT	50.25 42.615 51.405 42.72 ;
		RECT	50.25 43.11 51.405 43.2 ;
		RECT	51.21 43.2 51.405 43.61 ;
		RECT	50.25 43.3 51.11 43.51 ;
		RECT	50.25 43.61 51.405 43.705 ;
		RECT	51.21 43.705 51.405 44.095 ;
		RECT	50.25 44.095 51.405 44.2 ;
		RECT	50.25 44.59 51.405 44.685 ;
		RECT	50.25 45.075 51.405 45.18 ;
		RECT	50.25 45.57 51.405 45.655 ;
		RECT	51.21 45.655 51.405 46.655 ;
		RECT	50.25 46.055 51.11 46.265 ;
		RECT	50.25 46.38 51.1 46.57 ;
		RECT	51.21 47.19 51.405 47.495 ;
		RECT	50.25 47.245 51.11 47.435 ;
		RECT	50.25 48.03 51.405 48.13 ;
		RECT	50.25 48.52 51.405 48.62 ;
		RECT	50.25 49.01 51.405 49.115 ;
		RECT	50.25 49.505 51.405 49.605 ;
		RECT	50.25 49.995 51.405 50.1 ;
		RECT	51.21 50.635 51.405 50.935 ;
		RECT	50.25 50.69 51.11 50.88 ;
		RECT	51.21 51.47 51.405 52.47 ;
		RECT	50.25 51.495 51.11 51.685 ;
		RECT	50.25 51.83 51.11 52.04 ;
		RECT	50.25 52.47 51.405 52.555 ;
		RECT	50.25 52.945 51.405 53.05 ;
		RECT	50.25 53.44 51.405 53.545 ;
		RECT	50.25 53.935 51.405 54.025 ;
		RECT	51.21 54.025 51.405 54.435 ;
		RECT	50.25 54.435 51.405 54.515 ;
		RECT	51.21 54.515 51.405 54.925 ;
		RECT	50.25 54.615 51.11 54.825 ;
		RECT	50.25 54.925 51.405 55.02 ;
		RECT	50.25 55.41 51.405 55.51 ;
		RECT	50.25 55.9 51.405 56.005 ;
		RECT	50.25 56.395 51.405 56.485 ;
		RECT	50.25 56.895 51.405 56.985 ;
		RECT	50.25 57.375 51.405 57.48 ;
		RECT	50.25 57.87 51.405 57.97 ;
		RECT	50.25 58.36 51.405 58.465 ;
		RECT	51.21 58.465 51.405 58.855 ;
		RECT	50.25 58.565 51.11 58.755 ;
		RECT	50.25 58.855 51.405 58.955 ;
		RECT	50.25 59.345 51.405 59.445 ;
		RECT	50.25 59.835 51.405 59.94 ;
		RECT	50.25 60.33 51.405 60.43 ;
		RECT	50.25 60.82 51.405 60.925 ;
		RECT	50.25 61.315 51.405 61.415 ;
		RECT	50.25 61.805 51.405 61.905 ;
		RECT	50.65 62.295 51.405 62.39 ;
		RECT	51.21 62.39 51.405 62.8 ;
		RECT	50.25 62.49 51.11 62.7 ;
		RECT	50.25 62.8 51.405 62.89 ;
		RECT	50.25 63.28 51.405 63.375 ;
		RECT	51.03 63.375 51.405 63.785 ;
		RECT	50.98 63.785 51.405 63.875 ;
		RECT	50.98 64.265 51.405 64.355 ;
		RECT	50.25 64.765 51.405 64.825 ;
		RECT	50.25 65.215 51.405 65.35 ;
		RECT	50.25 65.74 51.405 65.81 ;
		RECT	51.21 66.2 51.405 66.69 ;
		RECT	50.25 66.2 51.11 66.35 ;
		RECT	50.25 66.45 51.11 66.64 ;
		RECT	51.21 66.87 51.405 67.215 ;
		RECT	50.25 66.925 51.11 67.115 ;
		RECT	50.25 67.215 51.405 67.32 ;
		RECT	50.25 68.2 51.405 68.305 ;
		RECT	51.21 68.695 51.405 69.045 ;
		RECT	50.25 68.705 51.11 68.915 ;
		RECT	50.25 69.045 51.405 69.155 ;
		RECT	50.25 69.885 51.405 71.285 ;
		RECT	14.49 29.15 23.73 29.34 ;
		RECT	14.49 29.825 23.73 29.925 ;
		RECT	14.49 30.805 23.73 30.91 ;
		RECT	14.49 31.01 23.73 31.2 ;
		RECT	14.49 31.485 23.73 31.675 ;
		RECT	14.49 31.775 14.74 31.93 ;
		RECT	14.8 31.78 23.73 31.93 ;
		RECT	14.49 32.32 23.73 32.385 ;
		RECT	14.49 32.775 23.73 32.88 ;
		RECT	14.49 33.27 23.73 33.37 ;
		RECT	14.49 34.25 23.73 34.355 ;
		RECT	14.49 34.745 23.73 34.845 ;
		RECT	14.49 35.235 23.73 35.34 ;
		RECT	14.49 35.44 23.73 35.63 ;
		RECT	14.49 35.73 23.73 35.83 ;
		RECT	14.49 36.22 23.73 36.325 ;
		RECT	14.49 36.715 23.73 36.815 ;
		RECT	14.49 37.205 23.73 37.305 ;
		RECT	14.49 37.695 23.73 37.8 ;
		RECT	14.49 38.19 23.73 38.29 ;
		RECT	14.49 38.68 23.73 38.78 ;
		RECT	14.49 39.17 23.73 39.275 ;
		RECT	14.49 39.375 23.73 39.565 ;
		RECT	14.49 39.665 23.73 39.765 ;
		RECT	14.49 40.155 23.73 40.26 ;
		RECT	14.49 40.65 23.73 40.75 ;
		RECT	14.49 41.14 23.73 41.23 ;
		RECT	14.49 41.64 23.73 41.735 ;
		RECT	14.49 42.125 23.73 42.225 ;
		RECT	14.49 42.615 23.73 42.72 ;
		RECT	14.49 43.11 23.73 43.2 ;
		RECT	14.49 43.3 23.73 43.51 ;
		RECT	14.49 43.61 23.73 43.705 ;
		RECT	14.49 44.095 23.73 44.2 ;
		RECT	14.49 44.59 23.73 44.685 ;
		RECT	14.49 45.075 23.73 45.18 ;
		RECT	14.49 45.57 23.73 45.655 ;
		RECT	14.49 46.045 14.7 46.28 ;
		RECT	14.8 46.055 23.73 46.265 ;
		RECT	14.49 46.38 23.73 46.57 ;
		RECT	14.49 47.245 23.73 47.435 ;
		RECT	14.49 48.03 23.73 48.13 ;
		RECT	14.49 48.52 23.73 48.62 ;
		RECT	14.49 49.01 23.73 49.115 ;
		RECT	14.49 49.505 23.73 49.605 ;
		RECT	14.49 49.995 23.73 50.1 ;
		RECT	14.49 50.69 23.73 50.88 ;
		RECT	14.49 51.495 23.73 51.685 ;
		RECT	14.49 51.785 14.7 52.08 ;
		RECT	14.8 51.83 23.73 52.04 ;
		RECT	14.49 52.47 23.73 52.555 ;
		RECT	14.49 52.945 23.73 53.05 ;
		RECT	14.49 53.44 23.73 53.545 ;
		RECT	14.49 53.935 23.73 54.025 ;
		RECT	14.49 54.435 23.73 54.515 ;
		RECT	14.49 54.615 23.73 54.825 ;
		RECT	14.49 54.925 23.73 55.02 ;
		RECT	14.49 55.41 23.73 55.51 ;
		RECT	14.49 55.9 23.73 56.005 ;
		RECT	14.49 56.395 23.73 56.485 ;
		RECT	14.49 56.895 23.73 56.985 ;
		RECT	14.49 57.375 23.73 57.48 ;
		RECT	14.49 57.87 23.73 57.97 ;
		RECT	14.49 58.36 23.73 58.465 ;
		RECT	14.49 58.565 23.73 58.755 ;
		RECT	14.49 58.855 23.73 58.955 ;
		RECT	14.49 59.345 23.73 59.445 ;
		RECT	14.49 59.835 23.73 59.94 ;
		RECT	14.49 60.33 23.73 60.43 ;
		RECT	14.49 60.82 23.73 60.925 ;
		RECT	14.49 61.315 23.73 61.415 ;
		RECT	14.49 61.805 23.73 61.905 ;
		RECT	14.49 62.49 23.73 62.7 ;
		RECT	14.49 62.8 23.73 62.89 ;
		RECT	14.49 63.28 23.73 63.375 ;
		RECT	14.49 63.79 23.73 63.86 ;
		RECT	14.49 64.28 23.73 64.35 ;
		RECT	14.49 64.765 23.73 64.825 ;
		RECT	14.49 65.215 23.73 65.35 ;
		RECT	14.49 65.74 23.73 65.81 ;
		RECT	14.49 66.2 14.74 66.35 ;
		RECT	14.8 66.2 23.73 66.35 ;
		RECT	14.49 66.45 23.73 66.64 ;
		RECT	14.49 66.925 23.73 67.115 ;
		RECT	14.49 67.215 23.73 67.32 ;
		RECT	14.49 68.2 23.73 68.305 ;
		RECT	14.49 68.705 23.73 68.915 ;
		RECT	23.73 29.15 24.27 29.34 ;
		RECT	23.73 29.825 24.27 29.925 ;
		RECT	23.73 30.805 24.27 30.91 ;
		RECT	23.73 31.01 24.27 31.2 ;
		RECT	23.73 31.485 24.27 31.675 ;
		RECT	23.73 31.78 24.27 31.93 ;
		RECT	23.73 32.32 24.27 32.385 ;
		RECT	23.73 32.775 24.27 32.88 ;
		RECT	23.73 33.27 24.27 33.37 ;
		RECT	23.73 34.25 24.27 34.355 ;
		RECT	23.73 34.745 24.27 34.845 ;
		RECT	23.73 35.235 24.27 35.34 ;
		RECT	23.73 35.44 24.27 35.63 ;
		RECT	23.73 35.73 24.27 35.83 ;
		RECT	23.73 36.22 24.27 36.325 ;
		RECT	23.73 36.715 24.27 36.815 ;
		RECT	23.73 37.205 24.27 37.305 ;
		RECT	23.73 37.695 24.27 37.8 ;
		RECT	23.73 38.19 24.27 38.29 ;
		RECT	23.73 38.68 24.27 38.78 ;
		RECT	23.73 39.17 24.27 39.275 ;
		RECT	23.73 39.375 24.27 39.565 ;
		RECT	23.73 39.665 24.27 39.765 ;
		RECT	23.73 40.155 24.27 40.26 ;
		RECT	23.73 40.65 24.27 40.75 ;
		RECT	23.73 41.14 24.27 41.23 ;
		RECT	23.73 41.64 24.27 41.735 ;
		RECT	23.73 42.125 24.27 42.225 ;
		RECT	23.73 42.615 24.27 42.72 ;
		RECT	23.73 43.11 24.27 43.2 ;
		RECT	23.73 43.3 24.27 43.51 ;
		RECT	23.73 43.61 24.27 43.705 ;
		RECT	23.73 44.095 24.27 44.2 ;
		RECT	23.73 44.59 24.27 44.685 ;
		RECT	23.73 45.075 24.27 45.18 ;
		RECT	23.73 45.57 24.27 45.655 ;
		RECT	23.73 46.055 24.27 46.265 ;
		RECT	23.73 46.38 24.27 46.57 ;
		RECT	23.73 47.245 24.27 47.435 ;
		RECT	23.73 48.03 24.27 48.13 ;
		RECT	23.73 48.52 24.27 48.62 ;
		RECT	23.73 49.01 24.27 49.115 ;
		RECT	23.73 49.505 24.27 49.605 ;
		RECT	23.73 49.995 24.27 50.1 ;
		RECT	23.73 50.69 24.27 50.88 ;
		RECT	23.73 51.495 24.27 51.685 ;
		RECT	23.73 51.83 24.27 52.04 ;
		RECT	23.73 52.47 24.27 52.555 ;
		RECT	23.73 52.945 24.27 53.05 ;
		RECT	23.73 53.44 24.27 53.545 ;
		RECT	23.73 53.935 24.27 54.025 ;
		RECT	23.73 54.435 24.27 54.515 ;
		RECT	23.73 54.615 24.27 54.825 ;
		RECT	23.73 54.925 24.27 55.02 ;
		RECT	23.73 55.41 24.27 55.51 ;
		RECT	23.73 55.9 24.27 56.005 ;
		RECT	23.73 56.395 24.27 56.485 ;
		RECT	23.73 56.895 24.27 56.985 ;
		RECT	23.73 57.375 24.27 57.48 ;
		RECT	23.73 57.87 24.27 57.97 ;
		RECT	23.73 58.36 24.27 58.465 ;
		RECT	23.73 58.565 24.27 58.755 ;
		RECT	23.73 58.855 24.27 58.955 ;
		RECT	23.73 59.345 24.27 59.445 ;
		RECT	23.73 59.835 24.27 59.94 ;
		RECT	23.73 60.33 24.27 60.43 ;
		RECT	23.73 60.82 24.27 60.925 ;
		RECT	23.73 61.315 24.27 61.415 ;
		RECT	23.73 61.805 24.27 61.905 ;
		RECT	23.73 62.49 24.27 62.7 ;
		RECT	23.73 62.8 24.27 62.89 ;
		RECT	23.73 63.28 24.27 63.375 ;
		RECT	23.73 63.79 24.27 63.86 ;
		RECT	23.73 64.28 24.27 64.35 ;
		RECT	23.73 64.765 24.27 64.825 ;
		RECT	23.73 65.215 24.27 65.35 ;
		RECT	23.73 65.74 24.27 65.81 ;
		RECT	23.73 66.2 24.27 66.35 ;
		RECT	23.73 66.45 24.27 66.64 ;
		RECT	23.73 66.925 24.27 67.115 ;
		RECT	23.73 67.215 24.27 67.32 ;
		RECT	23.73 68.2 24.27 68.305 ;
		RECT	23.73 68.705 24.27 68.915 ;
		RECT	24.27 29.15 24.81 29.34 ;
		RECT	24.27 29.825 24.81 29.925 ;
		RECT	24.27 30.805 24.81 30.91 ;
		RECT	24.27 31.01 24.81 31.2 ;
		RECT	24.27 31.485 24.81 31.675 ;
		RECT	24.27 31.78 24.81 31.93 ;
		RECT	24.27 32.32 24.81 32.385 ;
		RECT	24.27 32.775 24.81 32.88 ;
		RECT	24.27 33.27 24.81 33.37 ;
		RECT	24.27 34.25 24.81 34.355 ;
		RECT	24.27 34.745 24.81 34.845 ;
		RECT	24.27 35.235 24.81 35.34 ;
		RECT	24.27 35.44 24.81 35.63 ;
		RECT	24.27 35.73 24.81 35.83 ;
		RECT	24.27 36.22 24.81 36.325 ;
		RECT	24.27 36.715 24.81 36.815 ;
		RECT	24.27 37.205 24.81 37.305 ;
		RECT	24.27 37.695 24.81 37.8 ;
		RECT	24.27 38.19 24.81 38.29 ;
		RECT	24.27 38.68 24.81 38.78 ;
		RECT	24.27 39.17 24.81 39.275 ;
		RECT	24.27 39.375 24.81 39.565 ;
		RECT	24.27 39.665 24.81 39.765 ;
		RECT	24.27 40.155 24.81 40.26 ;
		RECT	24.27 40.65 24.81 40.75 ;
		RECT	24.27 41.14 24.81 41.23 ;
		RECT	24.27 41.64 24.81 41.735 ;
		RECT	24.27 42.125 24.81 42.225 ;
		RECT	24.27 42.615 24.81 42.72 ;
		RECT	24.27 43.11 24.81 43.2 ;
		RECT	24.27 43.3 24.81 43.51 ;
		RECT	24.27 43.61 24.81 43.705 ;
		RECT	24.27 44.095 24.81 44.2 ;
		RECT	24.27 44.59 24.81 44.685 ;
		RECT	24.27 45.075 24.81 45.18 ;
		RECT	24.27 45.57 24.81 45.655 ;
		RECT	24.27 46.055 24.81 46.265 ;
		RECT	24.27 46.38 24.81 46.57 ;
		RECT	24.27 47.245 24.81 47.435 ;
		RECT	24.27 48.03 24.81 48.13 ;
		RECT	24.27 48.52 24.81 48.62 ;
		RECT	24.27 49.01 24.81 49.115 ;
		RECT	24.27 49.505 24.81 49.605 ;
		RECT	24.27 49.995 24.81 50.1 ;
		RECT	24.27 50.69 24.81 50.88 ;
		RECT	24.27 51.495 24.81 51.685 ;
		RECT	24.27 51.83 24.81 52.04 ;
		RECT	24.27 52.47 24.81 52.555 ;
		RECT	24.27 52.945 24.81 53.05 ;
		RECT	24.27 53.44 24.81 53.545 ;
		RECT	24.27 53.935 24.81 54.025 ;
		RECT	24.27 54.435 24.81 54.515 ;
		RECT	24.27 54.615 24.81 54.825 ;
		RECT	24.27 54.925 24.81 55.02 ;
		RECT	24.27 55.41 24.81 55.51 ;
		RECT	24.27 55.9 24.81 56.005 ;
		RECT	24.27 56.395 24.81 56.485 ;
		RECT	24.27 56.895 24.81 56.985 ;
		RECT	24.27 57.375 24.81 57.48 ;
		RECT	24.27 57.87 24.81 57.97 ;
		RECT	24.27 58.36 24.81 58.465 ;
		RECT	24.27 58.565 24.81 58.755 ;
		RECT	24.27 58.855 24.81 58.955 ;
		RECT	24.27 59.345 24.81 59.445 ;
		RECT	24.27 59.835 24.81 59.94 ;
		RECT	24.27 60.33 24.81 60.43 ;
		RECT	24.27 60.82 24.81 60.925 ;
		RECT	24.27 61.315 24.81 61.415 ;
		RECT	24.27 61.805 24.81 61.905 ;
		RECT	24.27 62.49 24.81 62.7 ;
		RECT	24.27 62.8 24.81 62.89 ;
		RECT	24.27 63.28 24.81 63.375 ;
		RECT	24.27 63.79 24.81 63.86 ;
		RECT	24.27 64.28 24.81 64.35 ;
		RECT	24.27 64.765 24.81 64.825 ;
		RECT	24.27 65.215 24.81 65.35 ;
		RECT	24.27 65.74 24.81 65.81 ;
		RECT	24.27 66.2 24.81 66.35 ;
		RECT	24.27 66.45 24.81 66.64 ;
		RECT	24.27 66.925 24.81 67.115 ;
		RECT	24.27 67.215 24.81 67.32 ;
		RECT	24.27 68.2 24.81 68.305 ;
		RECT	24.27 68.705 24.81 68.915 ;
		RECT	24.81 29.15 25.35 29.34 ;
		RECT	24.81 29.825 25.35 29.925 ;
		RECT	24.81 30.805 25.35 30.91 ;
		RECT	24.81 31.01 25.35 31.2 ;
		RECT	24.81 31.485 25.35 31.675 ;
		RECT	24.81 31.78 25.35 31.93 ;
		RECT	24.81 32.32 25.35 32.385 ;
		RECT	24.81 32.775 25.35 32.88 ;
		RECT	24.81 33.27 25.35 33.37 ;
		RECT	24.81 34.25 25.35 34.355 ;
		RECT	24.81 34.745 25.35 34.845 ;
		RECT	24.81 35.235 25.35 35.34 ;
		RECT	24.81 35.44 25.35 35.63 ;
		RECT	24.81 35.73 25.35 35.83 ;
		RECT	24.81 36.22 25.35 36.325 ;
		RECT	24.81 36.715 25.35 36.815 ;
		RECT	24.81 37.205 25.35 37.305 ;
		RECT	24.81 37.695 25.35 37.8 ;
		RECT	24.81 38.19 25.35 38.29 ;
		RECT	24.81 38.68 25.35 38.78 ;
		RECT	24.81 39.17 25.35 39.275 ;
		RECT	24.81 39.375 25.35 39.565 ;
		RECT	24.81 39.665 25.35 39.765 ;
		RECT	24.81 40.155 25.35 40.26 ;
		RECT	24.81 40.65 25.35 40.75 ;
		RECT	24.81 41.14 25.35 41.23 ;
		RECT	24.81 41.64 25.35 41.735 ;
		RECT	24.81 42.125 25.35 42.225 ;
		RECT	24.81 42.615 25.35 42.72 ;
		RECT	24.81 43.11 25.35 43.2 ;
		RECT	24.81 43.3 25.35 43.51 ;
		RECT	24.81 43.61 25.35 43.705 ;
		RECT	24.81 44.095 25.35 44.2 ;
		RECT	24.81 44.59 25.35 44.685 ;
		RECT	24.81 45.075 25.35 45.18 ;
		RECT	24.81 45.57 25.35 45.655 ;
		RECT	24.81 46.055 25.35 46.265 ;
		RECT	24.81 46.38 25.35 46.57 ;
		RECT	24.81 47.245 25.35 47.435 ;
		RECT	24.81 48.03 25.35 48.13 ;
		RECT	24.81 48.52 25.35 48.62 ;
		RECT	24.81 49.01 25.35 49.115 ;
		RECT	24.81 49.505 25.35 49.605 ;
		RECT	24.81 49.995 25.35 50.1 ;
		RECT	24.81 50.69 25.35 50.88 ;
		RECT	24.81 51.495 25.35 51.685 ;
		RECT	24.81 51.83 25.35 52.04 ;
		RECT	24.81 52.47 25.35 52.555 ;
		RECT	24.81 52.945 25.35 53.05 ;
		RECT	24.81 53.44 25.35 53.545 ;
		RECT	24.81 53.935 25.35 54.025 ;
		RECT	24.81 54.435 25.35 54.515 ;
		RECT	24.81 54.615 25.35 54.825 ;
		RECT	24.81 54.925 25.35 55.02 ;
		RECT	24.81 55.41 25.35 55.51 ;
		RECT	24.81 55.9 25.35 56.005 ;
		RECT	24.81 56.395 25.35 56.485 ;
		RECT	24.81 56.895 25.35 56.985 ;
		RECT	24.81 57.375 25.35 57.48 ;
		RECT	24.81 57.87 25.35 57.97 ;
		RECT	24.81 58.36 25.35 58.465 ;
		RECT	24.81 58.565 25.35 58.755 ;
		RECT	24.81 58.855 25.35 58.955 ;
		RECT	24.81 59.345 25.35 59.445 ;
		RECT	24.81 59.835 25.35 59.94 ;
		RECT	24.81 60.33 25.35 60.43 ;
		RECT	24.81 60.82 25.35 60.925 ;
		RECT	24.81 61.315 25.35 61.415 ;
		RECT	24.81 61.805 25.35 61.905 ;
		RECT	24.81 62.49 25.35 62.7 ;
		RECT	24.81 62.8 25.35 62.89 ;
		RECT	24.81 63.28 25.35 63.375 ;
		RECT	24.81 63.79 25.35 63.86 ;
		RECT	24.81 64.28 25.35 64.35 ;
		RECT	24.81 64.765 25.35 64.825 ;
		RECT	24.81 65.215 25.35 65.35 ;
		RECT	24.81 65.74 25.35 65.81 ;
		RECT	24.81 66.2 25.35 66.35 ;
		RECT	24.81 66.45 25.35 66.64 ;
		RECT	24.81 66.925 25.35 67.115 ;
		RECT	24.81 67.215 25.35 67.32 ;
		RECT	24.81 68.2 25.35 68.305 ;
		RECT	24.81 68.705 25.35 68.915 ;
		RECT	25.35 29.15 25.89 29.34 ;
		RECT	25.35 29.825 25.89 29.925 ;
		RECT	25.35 30.805 25.89 30.91 ;
		RECT	25.35 31.01 25.89 31.2 ;
		RECT	25.35 31.485 25.89 31.675 ;
		RECT	25.35 31.78 25.89 31.93 ;
		RECT	25.35 32.32 25.89 32.385 ;
		RECT	25.35 32.775 25.89 32.88 ;
		RECT	25.35 33.27 25.89 33.37 ;
		RECT	25.35 34.25 25.89 34.355 ;
		RECT	25.35 34.745 25.89 34.845 ;
		RECT	25.35 35.235 25.89 35.34 ;
		RECT	25.35 35.44 25.89 35.63 ;
		RECT	25.35 35.73 25.89 35.83 ;
		RECT	25.35 36.22 25.89 36.325 ;
		RECT	25.35 36.715 25.89 36.815 ;
		RECT	25.35 37.205 25.89 37.305 ;
		RECT	25.35 37.695 25.89 37.8 ;
		RECT	25.35 38.19 25.89 38.29 ;
		RECT	25.35 38.68 25.89 38.78 ;
		RECT	25.35 39.17 25.89 39.275 ;
		RECT	25.35 39.375 25.89 39.565 ;
		RECT	25.35 39.665 25.89 39.765 ;
		RECT	25.35 40.155 25.89 40.26 ;
		RECT	25.35 40.65 25.89 40.75 ;
		RECT	25.35 41.14 25.89 41.23 ;
		RECT	25.35 41.64 25.89 41.735 ;
		RECT	25.35 42.125 25.89 42.225 ;
		RECT	25.35 42.615 25.89 42.72 ;
		RECT	25.35 43.11 25.89 43.2 ;
		RECT	25.35 43.3 25.89 43.51 ;
		RECT	25.35 43.61 25.89 43.705 ;
		RECT	25.35 44.095 25.89 44.2 ;
		RECT	25.35 44.59 25.89 44.685 ;
		RECT	25.35 45.075 25.89 45.18 ;
		RECT	25.35 45.57 25.89 45.655 ;
		RECT	25.35 46.055 25.89 46.265 ;
		RECT	25.35 46.38 25.89 46.57 ;
		RECT	25.35 47.245 25.89 47.435 ;
		RECT	25.35 48.03 25.89 48.13 ;
		RECT	25.35 48.52 25.89 48.62 ;
		RECT	25.35 49.01 25.89 49.115 ;
		RECT	25.35 49.505 25.89 49.605 ;
		RECT	25.35 49.995 25.89 50.1 ;
		RECT	25.35 50.69 25.89 50.88 ;
		RECT	25.35 51.495 25.89 51.685 ;
		RECT	25.35 51.83 25.89 52.04 ;
		RECT	25.35 52.47 25.89 52.555 ;
		RECT	25.35 52.945 25.89 53.05 ;
		RECT	25.35 53.44 25.89 53.545 ;
		RECT	25.35 53.935 25.89 54.025 ;
		RECT	25.35 54.435 25.89 54.515 ;
		RECT	25.35 54.615 25.89 54.825 ;
		RECT	25.35 54.925 25.89 55.02 ;
		RECT	25.35 55.41 25.89 55.51 ;
		RECT	25.35 55.9 25.89 56.005 ;
		RECT	25.35 56.395 25.89 56.485 ;
		RECT	25.35 56.895 25.89 56.985 ;
		RECT	25.35 57.375 25.89 57.48 ;
		RECT	25.35 57.87 25.89 57.97 ;
		RECT	25.35 58.36 25.89 58.465 ;
		RECT	25.35 58.565 25.89 58.755 ;
		RECT	25.35 58.855 25.89 58.955 ;
		RECT	25.35 59.345 25.89 59.445 ;
		RECT	25.35 59.835 25.89 59.94 ;
		RECT	25.35 60.33 25.89 60.43 ;
		RECT	25.35 60.82 25.89 60.925 ;
		RECT	25.35 61.315 25.89 61.415 ;
		RECT	25.35 61.805 25.89 61.905 ;
		RECT	25.35 62.49 25.89 62.7 ;
		RECT	25.35 62.8 25.89 62.89 ;
		RECT	25.35 63.28 25.89 63.375 ;
		RECT	25.35 63.79 25.89 63.86 ;
		RECT	25.35 64.28 25.89 64.35 ;
		RECT	25.35 64.765 25.89 64.825 ;
		RECT	25.35 65.215 25.89 65.35 ;
		RECT	25.35 65.74 25.89 65.81 ;
		RECT	25.35 66.2 25.89 66.35 ;
		RECT	25.35 66.45 25.89 66.64 ;
		RECT	25.35 66.925 25.89 67.115 ;
		RECT	25.35 67.215 25.89 67.32 ;
		RECT	25.35 68.2 25.89 68.305 ;
		RECT	25.35 68.705 25.89 68.915 ;
		RECT	25.89 29.15 26.43 29.34 ;
		RECT	25.89 29.825 26.43 29.925 ;
		RECT	25.89 30.805 26.43 30.91 ;
		RECT	25.89 31.01 26.43 31.2 ;
		RECT	25.89 31.485 26.43 31.675 ;
		RECT	25.89 31.78 26.43 31.93 ;
		RECT	25.89 32.32 26.43 32.385 ;
		RECT	25.89 32.775 26.43 32.88 ;
		RECT	25.89 33.27 26.43 33.37 ;
		RECT	25.89 34.25 26.43 34.355 ;
		RECT	25.89 34.745 26.43 34.845 ;
		RECT	25.89 35.235 26.43 35.34 ;
		RECT	25.89 35.44 26.43 35.63 ;
		RECT	25.89 35.73 26.43 35.83 ;
		RECT	25.89 36.22 26.43 36.325 ;
		RECT	25.89 36.715 26.43 36.815 ;
		RECT	25.89 37.205 26.43 37.305 ;
		RECT	25.89 37.695 26.43 37.8 ;
		RECT	25.89 38.19 26.43 38.29 ;
		RECT	25.89 38.68 26.43 38.78 ;
		RECT	25.89 39.17 26.43 39.275 ;
		RECT	25.89 39.375 26.43 39.565 ;
		RECT	25.89 39.665 26.43 39.765 ;
		RECT	25.89 40.155 26.43 40.26 ;
		RECT	25.89 40.65 26.43 40.75 ;
		RECT	25.89 41.14 26.43 41.23 ;
		RECT	25.89 41.64 26.43 41.735 ;
		RECT	25.89 42.125 26.43 42.225 ;
		RECT	25.89 42.615 26.43 42.72 ;
		RECT	25.89 43.11 26.43 43.2 ;
		RECT	25.89 43.3 26.43 43.51 ;
		RECT	25.89 43.61 26.43 43.705 ;
		RECT	25.89 44.095 26.43 44.2 ;
		RECT	25.89 44.59 26.43 44.685 ;
		RECT	25.89 45.075 26.43 45.18 ;
		RECT	25.89 45.57 26.43 45.655 ;
		RECT	25.89 46.055 26.43 46.265 ;
		RECT	25.89 46.38 26.43 46.57 ;
		RECT	25.89 47.245 26.43 47.435 ;
		RECT	25.89 48.03 26.43 48.13 ;
		RECT	25.89 48.52 26.43 48.62 ;
		RECT	25.89 49.01 26.43 49.115 ;
		RECT	25.89 49.505 26.43 49.605 ;
		RECT	25.89 49.995 26.43 50.1 ;
		RECT	25.89 50.69 26.43 50.88 ;
		RECT	25.89 51.495 26.43 51.685 ;
		RECT	25.89 51.83 26.43 52.04 ;
		RECT	25.89 52.47 26.43 52.555 ;
		RECT	25.89 52.945 26.43 53.05 ;
		RECT	25.89 53.44 26.43 53.545 ;
		RECT	25.89 53.935 26.43 54.025 ;
		RECT	25.89 54.435 26.43 54.515 ;
		RECT	25.89 54.615 26.43 54.825 ;
		RECT	25.89 54.925 26.43 55.02 ;
		RECT	25.89 55.41 26.43 55.51 ;
		RECT	25.89 55.9 26.43 56.005 ;
		RECT	25.89 56.395 26.43 56.485 ;
		RECT	25.89 56.895 26.43 56.985 ;
		RECT	25.89 57.375 26.43 57.48 ;
		RECT	25.89 57.87 26.43 57.97 ;
		RECT	25.89 58.36 26.43 58.465 ;
		RECT	25.89 58.565 26.43 58.755 ;
		RECT	25.89 58.855 26.43 58.955 ;
		RECT	25.89 59.345 26.43 59.445 ;
		RECT	25.89 59.835 26.43 59.94 ;
		RECT	25.89 60.33 26.43 60.43 ;
		RECT	25.89 60.82 26.43 60.925 ;
		RECT	25.89 61.315 26.43 61.415 ;
		RECT	25.89 61.805 26.43 61.905 ;
		RECT	25.89 62.49 26.43 62.7 ;
		RECT	25.89 62.8 26.43 62.89 ;
		RECT	25.89 63.28 26.43 63.375 ;
		RECT	25.89 63.79 26.43 63.86 ;
		RECT	25.89 64.28 26.43 64.35 ;
		RECT	25.89 64.765 26.43 64.825 ;
		RECT	25.89 65.215 26.43 65.35 ;
		RECT	25.89 65.74 26.43 65.81 ;
		RECT	25.89 66.2 26.43 66.35 ;
		RECT	25.89 66.45 26.43 66.64 ;
		RECT	25.89 66.925 26.43 67.115 ;
		RECT	25.89 67.215 26.43 67.32 ;
		RECT	25.89 68.2 26.43 68.305 ;
		RECT	25.89 68.705 26.43 68.915 ;
		RECT	26.43 29.15 26.97 29.34 ;
		RECT	26.43 29.825 26.97 29.925 ;
		RECT	26.43 30.805 26.97 30.91 ;
		RECT	26.43 31.01 26.97 31.2 ;
		RECT	26.43 31.485 26.97 31.675 ;
		RECT	26.43 31.78 26.97 31.93 ;
		RECT	26.43 32.32 26.97 32.385 ;
		RECT	26.43 32.775 26.97 32.88 ;
		RECT	26.43 33.27 26.97 33.37 ;
		RECT	26.43 34.25 26.97 34.355 ;
		RECT	26.43 34.745 26.97 34.845 ;
		RECT	26.43 35.235 26.97 35.34 ;
		RECT	26.43 35.44 26.97 35.63 ;
		RECT	26.43 35.73 26.97 35.83 ;
		RECT	26.43 36.22 26.97 36.325 ;
		RECT	26.43 36.715 26.97 36.815 ;
		RECT	26.43 37.205 26.97 37.305 ;
		RECT	26.43 37.695 26.97 37.8 ;
		RECT	26.43 38.19 26.97 38.29 ;
		RECT	26.43 38.68 26.97 38.78 ;
		RECT	26.43 39.17 26.97 39.275 ;
		RECT	26.43 39.375 26.97 39.565 ;
		RECT	26.43 39.665 26.97 39.765 ;
		RECT	26.43 40.155 26.97 40.26 ;
		RECT	26.43 40.65 26.97 40.75 ;
		RECT	26.43 41.14 26.97 41.23 ;
		RECT	26.43 41.64 26.97 41.735 ;
		RECT	26.43 42.125 26.97 42.225 ;
		RECT	26.43 42.615 26.97 42.72 ;
		RECT	26.43 43.11 26.97 43.2 ;
		RECT	26.43 43.3 26.97 43.51 ;
		RECT	26.43 43.61 26.97 43.705 ;
		RECT	26.43 44.095 26.97 44.2 ;
		RECT	26.43 44.59 26.97 44.685 ;
		RECT	26.43 45.075 26.97 45.18 ;
		RECT	26.43 45.57 26.97 45.655 ;
		RECT	26.43 46.055 26.97 46.265 ;
		RECT	26.43 46.38 26.97 46.57 ;
		RECT	26.43 47.245 26.97 47.435 ;
		RECT	26.43 48.03 26.97 48.13 ;
		RECT	26.43 48.52 26.97 48.62 ;
		RECT	26.43 49.01 26.97 49.115 ;
		RECT	26.43 49.505 26.97 49.605 ;
		RECT	26.43 49.995 26.97 50.1 ;
		RECT	26.43 50.69 26.97 50.88 ;
		RECT	26.43 51.495 26.97 51.685 ;
		RECT	26.43 51.83 26.97 52.04 ;
		RECT	26.43 52.47 26.97 52.555 ;
		RECT	26.43 52.945 26.97 53.05 ;
		RECT	26.43 53.44 26.97 53.545 ;
		RECT	26.43 53.935 26.97 54.025 ;
		RECT	26.43 54.435 26.97 54.515 ;
		RECT	26.43 54.615 26.97 54.825 ;
		RECT	26.43 54.925 26.97 55.02 ;
		RECT	26.43 55.41 26.97 55.51 ;
		RECT	26.43 55.9 26.97 56.005 ;
		RECT	26.43 56.395 26.97 56.485 ;
		RECT	26.43 56.895 26.97 56.985 ;
		RECT	26.43 57.375 26.97 57.48 ;
		RECT	26.43 57.87 26.97 57.97 ;
		RECT	26.43 58.36 26.97 58.465 ;
		RECT	26.43 58.565 26.97 58.755 ;
		RECT	26.43 58.855 26.97 58.955 ;
		RECT	26.43 59.345 26.97 59.445 ;
		RECT	26.43 59.835 26.97 59.94 ;
		RECT	26.43 60.33 26.97 60.43 ;
		RECT	26.43 60.82 26.97 60.925 ;
		RECT	26.43 61.315 26.97 61.415 ;
		RECT	26.43 61.805 26.97 61.905 ;
		RECT	26.43 62.49 26.97 62.7 ;
		RECT	26.43 62.8 26.97 62.89 ;
		RECT	26.43 63.28 26.97 63.375 ;
		RECT	26.43 63.79 26.97 63.86 ;
		RECT	26.43 64.28 26.97 64.35 ;
		RECT	26.43 64.765 26.97 64.825 ;
		RECT	26.43 65.215 26.97 65.35 ;
		RECT	26.43 65.74 26.97 65.81 ;
		RECT	26.43 66.2 26.97 66.35 ;
		RECT	26.43 66.45 26.97 66.64 ;
		RECT	26.43 66.925 26.97 67.115 ;
		RECT	26.43 67.215 26.97 67.32 ;
		RECT	26.43 68.2 26.97 68.305 ;
		RECT	26.43 68.705 26.97 68.915 ;
		RECT	26.97 29.15 27.51 29.34 ;
		RECT	26.97 29.825 27.51 29.925 ;
		RECT	26.97 30.805 27.51 30.91 ;
		RECT	26.97 31.01 27.51 31.2 ;
		RECT	26.97 31.485 27.51 31.675 ;
		RECT	26.97 31.78 27.51 31.93 ;
		RECT	26.97 32.32 27.51 32.385 ;
		RECT	26.97 32.775 27.51 32.88 ;
		RECT	26.97 33.27 27.51 33.37 ;
		RECT	26.97 34.25 27.51 34.355 ;
		RECT	26.97 34.745 27.51 34.845 ;
		RECT	26.97 35.235 27.51 35.34 ;
		RECT	26.97 35.44 27.51 35.63 ;
		RECT	26.97 35.73 27.51 35.83 ;
		RECT	26.97 36.22 27.51 36.325 ;
		RECT	26.97 36.715 27.51 36.815 ;
		RECT	26.97 37.205 27.51 37.305 ;
		RECT	26.97 37.695 27.51 37.8 ;
		RECT	26.97 38.19 27.51 38.29 ;
		RECT	26.97 38.68 27.51 38.78 ;
		RECT	26.97 39.17 27.51 39.275 ;
		RECT	26.97 39.375 27.51 39.565 ;
		RECT	26.97 39.665 27.51 39.765 ;
		RECT	26.97 40.155 27.51 40.26 ;
		RECT	26.97 40.65 27.51 40.75 ;
		RECT	26.97 41.14 27.51 41.23 ;
		RECT	26.97 41.64 27.51 41.735 ;
		RECT	26.97 42.125 27.51 42.225 ;
		RECT	26.97 42.615 27.51 42.72 ;
		RECT	26.97 43.11 27.51 43.2 ;
		RECT	26.97 43.3 27.51 43.51 ;
		RECT	26.97 43.61 27.51 43.705 ;
		RECT	26.97 44.095 27.51 44.2 ;
		RECT	26.97 44.59 27.51 44.685 ;
		RECT	26.97 45.075 27.51 45.18 ;
		RECT	26.97 45.57 27.51 45.655 ;
		RECT	26.97 46.055 27.51 46.265 ;
		RECT	26.97 46.38 27.51 46.57 ;
		RECT	26.97 47.245 27.51 47.435 ;
		RECT	26.97 48.03 27.51 48.13 ;
		RECT	26.97 48.52 27.51 48.62 ;
		RECT	26.97 49.01 27.51 49.115 ;
		RECT	26.97 49.505 27.51 49.605 ;
		RECT	26.97 49.995 27.51 50.1 ;
		RECT	26.97 50.69 27.51 50.88 ;
		RECT	26.97 51.495 27.51 51.685 ;
		RECT	26.97 51.83 27.51 52.04 ;
		RECT	26.97 52.47 27.51 52.555 ;
		RECT	26.97 52.945 27.51 53.05 ;
		RECT	26.97 53.44 27.51 53.545 ;
		RECT	26.97 53.935 27.51 54.025 ;
		RECT	26.97 54.435 27.51 54.515 ;
		RECT	26.97 54.615 27.51 54.825 ;
		RECT	26.97 54.925 27.51 55.02 ;
		RECT	26.97 55.41 27.51 55.51 ;
		RECT	26.97 55.9 27.51 56.005 ;
		RECT	26.97 56.395 27.51 56.485 ;
		RECT	26.97 56.895 27.51 56.985 ;
		RECT	26.97 57.375 27.51 57.48 ;
		RECT	26.97 57.87 27.51 57.97 ;
		RECT	26.97 58.36 27.51 58.465 ;
		RECT	26.97 58.565 27.51 58.755 ;
		RECT	26.97 58.855 27.51 58.955 ;
		RECT	26.97 59.345 27.51 59.445 ;
		RECT	26.97 59.835 27.51 59.94 ;
		RECT	26.97 60.33 27.51 60.43 ;
		RECT	26.97 60.82 27.51 60.925 ;
		RECT	26.97 61.315 27.51 61.415 ;
		RECT	26.97 61.805 27.51 61.905 ;
		RECT	26.97 62.49 27.51 62.7 ;
		RECT	26.97 62.8 27.51 62.89 ;
		RECT	26.97 63.28 27.51 63.375 ;
		RECT	26.97 63.79 27.51 63.86 ;
		RECT	26.97 64.28 27.51 64.35 ;
		RECT	26.97 64.765 27.51 64.825 ;
		RECT	26.97 65.215 27.51 65.35 ;
		RECT	26.97 65.74 27.51 65.81 ;
		RECT	26.97 66.2 27.51 66.35 ;
		RECT	26.97 66.45 27.51 66.64 ;
		RECT	26.97 66.925 27.51 67.115 ;
		RECT	26.97 67.215 27.51 67.32 ;
		RECT	26.97 68.2 27.51 68.305 ;
		RECT	26.97 68.705 27.51 68.915 ;
		RECT	27.51 29.15 28.05 29.34 ;
		RECT	27.51 29.825 28.05 29.925 ;
		RECT	27.51 30.805 28.05 30.91 ;
		RECT	27.51 31.01 28.05 31.2 ;
		RECT	27.51 31.485 28.05 31.675 ;
		RECT	27.51 31.78 28.05 31.93 ;
		RECT	27.51 32.32 28.05 32.385 ;
		RECT	27.51 32.775 28.05 32.88 ;
		RECT	27.51 33.27 28.05 33.37 ;
		RECT	27.51 34.25 28.05 34.355 ;
		RECT	27.51 34.745 28.05 34.845 ;
		RECT	27.51 35.235 28.05 35.34 ;
		RECT	27.51 35.44 28.05 35.63 ;
		RECT	27.51 35.73 28.05 35.83 ;
		RECT	27.51 36.22 28.05 36.325 ;
		RECT	27.51 36.715 28.05 36.815 ;
		RECT	27.51 37.205 28.05 37.305 ;
		RECT	27.51 37.695 28.05 37.8 ;
		RECT	27.51 38.19 28.05 38.29 ;
		RECT	27.51 38.68 28.05 38.78 ;
		RECT	27.51 39.17 28.05 39.275 ;
		RECT	27.51 39.375 28.05 39.565 ;
		RECT	27.51 39.665 28.05 39.765 ;
		RECT	27.51 40.155 28.05 40.26 ;
		RECT	27.51 40.65 28.05 40.75 ;
		RECT	27.51 41.14 28.05 41.23 ;
		RECT	27.51 41.64 28.05 41.735 ;
		RECT	27.51 42.125 28.05 42.225 ;
		RECT	27.51 42.615 28.05 42.72 ;
		RECT	27.51 43.11 28.05 43.2 ;
		RECT	27.51 43.3 28.05 43.51 ;
		RECT	27.51 43.61 28.05 43.705 ;
		RECT	27.51 44.095 28.05 44.2 ;
		RECT	27.51 44.59 28.05 44.685 ;
		RECT	27.51 45.075 28.05 45.18 ;
		RECT	27.51 45.57 28.05 45.655 ;
		RECT	27.51 46.055 28.05 46.265 ;
		RECT	27.51 46.38 28.05 46.57 ;
		RECT	27.51 47.245 28.05 47.435 ;
		RECT	27.51 48.03 28.05 48.13 ;
		RECT	27.51 48.52 28.05 48.62 ;
		RECT	27.51 49.01 28.05 49.115 ;
		RECT	27.51 49.505 28.05 49.605 ;
		RECT	27.51 49.995 28.05 50.1 ;
		RECT	27.51 50.69 28.05 50.88 ;
		RECT	27.51 51.495 28.05 51.685 ;
		RECT	27.51 51.83 28.05 52.04 ;
		RECT	27.51 52.47 28.05 52.555 ;
		RECT	27.51 52.945 28.05 53.05 ;
		RECT	27.51 53.44 28.05 53.545 ;
		RECT	27.51 53.935 28.05 54.025 ;
		RECT	27.51 54.435 28.05 54.515 ;
		RECT	27.51 54.615 28.05 54.825 ;
		RECT	27.51 54.925 28.05 55.02 ;
		RECT	27.51 55.41 28.05 55.51 ;
		RECT	27.51 55.9 28.05 56.005 ;
		RECT	27.51 56.395 28.05 56.485 ;
		RECT	27.51 56.895 28.05 56.985 ;
		RECT	27.51 57.375 28.05 57.48 ;
		RECT	27.51 57.87 28.05 57.97 ;
		RECT	27.51 58.36 28.05 58.465 ;
		RECT	27.51 58.565 28.05 58.755 ;
		RECT	27.51 58.855 28.05 58.955 ;
		RECT	27.51 59.345 28.05 59.445 ;
		RECT	27.51 59.835 28.05 59.94 ;
		RECT	27.51 60.33 28.05 60.43 ;
		RECT	27.51 60.82 28.05 60.925 ;
		RECT	27.51 61.315 28.05 61.415 ;
		RECT	27.51 61.805 28.05 61.905 ;
		RECT	27.51 62.49 28.05 62.7 ;
		RECT	27.51 62.8 28.05 62.89 ;
		RECT	27.51 63.28 28.05 63.375 ;
		RECT	27.51 63.79 28.05 63.86 ;
		RECT	27.51 64.28 28.05 64.35 ;
		RECT	27.51 64.765 28.05 64.825 ;
		RECT	27.51 65.215 28.05 65.35 ;
		RECT	27.51 65.74 28.05 65.81 ;
		RECT	27.51 66.2 28.05 66.35 ;
		RECT	27.51 66.45 28.05 66.64 ;
		RECT	27.51 66.925 28.05 67.115 ;
		RECT	27.51 67.215 28.05 67.32 ;
		RECT	27.51 68.2 28.05 68.305 ;
		RECT	27.51 68.705 28.05 68.915 ;
		RECT	28.05 29.15 28.59 29.34 ;
		RECT	28.05 29.825 28.59 29.925 ;
		RECT	28.05 30.805 28.59 30.91 ;
		RECT	28.05 31.01 28.59 31.2 ;
		RECT	28.05 31.485 28.59 31.675 ;
		RECT	28.05 31.78 28.59 31.93 ;
		RECT	28.05 32.32 28.59 32.385 ;
		RECT	28.05 32.775 28.59 32.88 ;
		RECT	28.05 33.27 28.59 33.37 ;
		RECT	28.05 34.25 28.59 34.355 ;
		RECT	28.05 34.745 28.59 34.845 ;
		RECT	28.05 35.235 28.59 35.34 ;
		RECT	28.05 35.44 28.59 35.63 ;
		RECT	28.05 35.73 28.59 35.83 ;
		RECT	28.05 36.22 28.59 36.325 ;
		RECT	28.05 36.715 28.59 36.815 ;
		RECT	28.05 37.205 28.59 37.305 ;
		RECT	28.05 37.695 28.59 37.8 ;
		RECT	28.05 38.19 28.59 38.29 ;
		RECT	28.05 38.68 28.59 38.78 ;
		RECT	28.05 39.17 28.59 39.275 ;
		RECT	28.05 39.375 28.59 39.565 ;
		RECT	28.05 39.665 28.59 39.765 ;
		RECT	28.05 40.155 28.59 40.26 ;
		RECT	28.05 40.65 28.59 40.75 ;
		RECT	28.05 41.14 28.59 41.23 ;
		RECT	28.05 41.64 28.59 41.735 ;
		RECT	28.05 42.125 28.59 42.225 ;
		RECT	28.05 42.615 28.59 42.72 ;
		RECT	28.05 43.11 28.59 43.2 ;
		RECT	28.05 43.3 28.59 43.51 ;
		RECT	28.05 43.61 28.59 43.705 ;
		RECT	28.05 44.095 28.59 44.2 ;
		RECT	28.05 44.59 28.59 44.685 ;
		RECT	28.05 45.075 28.59 45.18 ;
		RECT	28.05 45.57 28.59 45.655 ;
		RECT	28.05 46.055 28.59 46.265 ;
		RECT	28.05 46.38 28.59 46.57 ;
		RECT	28.05 47.245 28.59 47.435 ;
		RECT	28.05 48.03 28.59 48.13 ;
		RECT	28.05 48.52 28.59 48.62 ;
		RECT	28.05 49.01 28.59 49.115 ;
		RECT	28.05 49.505 28.59 49.605 ;
		RECT	28.05 49.995 28.59 50.1 ;
		RECT	28.05 50.69 28.59 50.88 ;
		RECT	28.05 51.495 28.59 51.685 ;
		RECT	28.05 51.83 28.59 52.04 ;
		RECT	28.05 52.47 28.59 52.555 ;
		RECT	28.05 52.945 28.59 53.05 ;
		RECT	28.05 53.44 28.59 53.545 ;
		RECT	28.05 53.935 28.59 54.025 ;
		RECT	28.05 54.435 28.59 54.515 ;
		RECT	28.05 54.615 28.59 54.825 ;
		RECT	28.05 54.925 28.59 55.02 ;
		RECT	28.05 55.41 28.59 55.51 ;
		RECT	28.05 55.9 28.59 56.005 ;
		RECT	28.05 56.395 28.59 56.485 ;
		RECT	28.05 56.895 28.59 56.985 ;
		RECT	28.05 57.375 28.59 57.48 ;
		RECT	28.05 57.87 28.59 57.97 ;
		RECT	28.05 58.36 28.59 58.465 ;
		RECT	28.05 58.565 28.59 58.755 ;
		RECT	28.05 58.855 28.59 58.955 ;
		RECT	28.05 59.345 28.59 59.445 ;
		RECT	28.05 59.835 28.59 59.94 ;
		RECT	28.05 60.33 28.59 60.43 ;
		RECT	28.05 60.82 28.59 60.925 ;
		RECT	28.05 61.315 28.59 61.415 ;
		RECT	28.05 61.805 28.59 61.905 ;
		RECT	28.05 62.49 28.59 62.7 ;
		RECT	28.05 62.8 28.59 62.89 ;
		RECT	28.05 63.28 28.59 63.375 ;
		RECT	28.05 63.79 28.59 63.86 ;
		RECT	28.05 64.28 28.59 64.35 ;
		RECT	28.05 64.765 28.59 64.825 ;
		RECT	28.05 65.215 28.59 65.35 ;
		RECT	28.05 65.74 28.59 65.81 ;
		RECT	28.05 66.2 28.59 66.35 ;
		RECT	28.05 66.45 28.59 66.64 ;
		RECT	28.05 66.925 28.59 67.115 ;
		RECT	28.05 67.215 28.59 67.32 ;
		RECT	28.05 68.2 28.59 68.305 ;
		RECT	28.05 68.705 28.59 68.915 ;
		RECT	28.59 29.15 29.13 29.34 ;
		RECT	28.59 29.825 29.13 29.925 ;
		RECT	28.59 30.805 29.13 30.91 ;
		RECT	28.59 31.01 29.13 31.2 ;
		RECT	28.59 31.485 29.13 31.675 ;
		RECT	28.59 31.78 29.13 31.93 ;
		RECT	28.59 32.32 29.13 32.385 ;
		RECT	28.59 32.775 29.13 32.88 ;
		RECT	28.59 33.27 29.13 33.37 ;
		RECT	28.59 34.25 29.13 34.355 ;
		RECT	28.59 34.745 29.13 34.845 ;
		RECT	28.59 35.235 29.13 35.34 ;
		RECT	28.59 35.44 29.13 35.63 ;
		RECT	28.59 35.73 29.13 35.83 ;
		RECT	28.59 36.22 29.13 36.325 ;
		RECT	28.59 36.715 29.13 36.815 ;
		RECT	28.59 37.205 29.13 37.305 ;
		RECT	28.59 37.695 29.13 37.8 ;
		RECT	28.59 38.19 29.13 38.29 ;
		RECT	28.59 38.68 29.13 38.78 ;
		RECT	28.59 39.17 29.13 39.275 ;
		RECT	28.59 39.375 29.13 39.565 ;
		RECT	28.59 39.665 29.13 39.765 ;
		RECT	28.59 40.155 29.13 40.26 ;
		RECT	28.59 40.65 29.13 40.75 ;
		RECT	28.59 41.14 29.13 41.23 ;
		RECT	28.59 41.64 29.13 41.735 ;
		RECT	28.59 42.125 29.13 42.225 ;
		RECT	28.59 42.615 29.13 42.72 ;
		RECT	28.59 43.11 29.13 43.2 ;
		RECT	28.59 43.3 29.13 43.51 ;
		RECT	28.59 43.61 29.13 43.705 ;
		RECT	28.59 44.095 29.13 44.2 ;
		RECT	28.59 44.59 29.13 44.685 ;
		RECT	28.59 45.075 29.13 45.18 ;
		RECT	28.59 45.57 29.13 45.655 ;
		RECT	28.59 46.055 29.13 46.265 ;
		RECT	28.59 46.38 29.13 46.57 ;
		RECT	28.59 47.245 29.13 47.435 ;
		RECT	28.59 48.03 29.13 48.13 ;
		RECT	28.59 48.52 29.13 48.62 ;
		RECT	28.59 49.01 29.13 49.115 ;
		RECT	28.59 49.505 29.13 49.605 ;
		RECT	28.59 49.995 29.13 50.1 ;
		RECT	28.59 50.69 29.13 50.88 ;
		RECT	28.59 51.495 29.13 51.685 ;
		RECT	28.59 51.83 29.13 52.04 ;
		RECT	28.59 52.47 29.13 52.555 ;
		RECT	28.59 52.945 29.13 53.05 ;
		RECT	28.59 53.44 29.13 53.545 ;
		RECT	28.59 53.935 29.13 54.025 ;
		RECT	28.59 54.435 29.13 54.515 ;
		RECT	28.59 54.615 29.13 54.825 ;
		RECT	28.59 54.925 29.13 55.02 ;
		RECT	28.59 55.41 29.13 55.51 ;
		RECT	28.59 55.9 29.13 56.005 ;
		RECT	28.59 56.395 29.13 56.485 ;
		RECT	28.59 56.895 29.13 56.985 ;
		RECT	28.59 57.375 29.13 57.48 ;
		RECT	28.59 57.87 29.13 57.97 ;
		RECT	28.59 58.36 29.13 58.465 ;
		RECT	28.59 58.565 29.13 58.755 ;
		RECT	28.59 58.855 29.13 58.955 ;
		RECT	28.59 59.345 29.13 59.445 ;
		RECT	28.59 59.835 29.13 59.94 ;
		RECT	28.59 60.33 29.13 60.43 ;
		RECT	28.59 60.82 29.13 60.925 ;
		RECT	28.59 61.315 29.13 61.415 ;
		RECT	28.59 61.805 29.13 61.905 ;
		RECT	28.59 62.49 29.13 62.7 ;
		RECT	28.59 62.8 29.13 62.89 ;
		RECT	28.59 63.28 29.13 63.375 ;
		RECT	28.59 63.79 29.13 63.86 ;
		RECT	28.59 64.28 29.13 64.35 ;
		RECT	28.59 64.765 29.13 64.825 ;
		RECT	28.59 65.215 29.13 65.35 ;
		RECT	28.59 65.74 29.13 65.81 ;
		RECT	28.59 66.2 29.13 66.35 ;
		RECT	28.59 66.45 29.13 66.64 ;
		RECT	28.59 66.925 29.13 67.115 ;
		RECT	28.59 67.215 29.13 67.32 ;
		RECT	28.59 68.2 29.13 68.305 ;
		RECT	28.59 68.705 29.13 68.915 ;
		RECT	29.13 29.15 29.67 29.34 ;
		RECT	29.13 29.825 29.67 29.925 ;
		RECT	29.13 30.805 29.67 30.91 ;
		RECT	29.13 31.01 29.67 31.2 ;
		RECT	29.13 31.485 29.67 31.675 ;
		RECT	29.13 31.78 29.67 31.93 ;
		RECT	29.13 32.32 29.67 32.385 ;
		RECT	29.13 32.775 29.67 32.88 ;
		RECT	29.13 33.27 29.67 33.37 ;
		RECT	29.13 34.25 29.67 34.355 ;
		RECT	29.13 34.745 29.67 34.845 ;
		RECT	29.13 35.235 29.67 35.34 ;
		RECT	29.13 35.44 29.67 35.63 ;
		RECT	29.13 35.73 29.67 35.83 ;
		RECT	29.13 36.22 29.67 36.325 ;
		RECT	29.13 36.715 29.67 36.815 ;
		RECT	29.13 37.205 29.67 37.305 ;
		RECT	29.13 37.695 29.67 37.8 ;
		RECT	29.13 38.19 29.67 38.29 ;
		RECT	29.13 38.68 29.67 38.78 ;
		RECT	29.13 39.17 29.67 39.275 ;
		RECT	29.13 39.375 29.67 39.565 ;
		RECT	29.13 39.665 29.67 39.765 ;
		RECT	29.13 40.155 29.67 40.26 ;
		RECT	29.13 40.65 29.67 40.75 ;
		RECT	29.13 41.14 29.67 41.23 ;
		RECT	29.13 41.64 29.67 41.735 ;
		RECT	29.13 42.125 29.67 42.225 ;
		RECT	29.13 42.615 29.67 42.72 ;
		RECT	29.13 43.11 29.67 43.2 ;
		RECT	29.13 43.3 29.67 43.51 ;
		RECT	29.13 43.61 29.67 43.705 ;
		RECT	29.13 44.095 29.67 44.2 ;
		RECT	29.13 44.59 29.67 44.685 ;
		RECT	29.13 45.075 29.67 45.18 ;
		RECT	29.13 45.57 29.67 45.655 ;
		RECT	29.13 46.055 29.67 46.265 ;
		RECT	29.13 46.38 29.67 46.57 ;
		RECT	29.13 47.245 29.67 47.435 ;
		RECT	29.13 48.03 29.67 48.13 ;
		RECT	29.13 48.52 29.67 48.62 ;
		RECT	29.13 49.01 29.67 49.115 ;
		RECT	29.13 49.505 29.67 49.605 ;
		RECT	29.13 49.995 29.67 50.1 ;
		RECT	29.13 50.69 29.67 50.88 ;
		RECT	29.13 51.495 29.67 51.685 ;
		RECT	29.13 51.83 29.67 52.04 ;
		RECT	29.13 52.47 29.67 52.555 ;
		RECT	29.13 52.945 29.67 53.05 ;
		RECT	29.13 53.44 29.67 53.545 ;
		RECT	29.13 53.935 29.67 54.025 ;
		RECT	29.13 54.435 29.67 54.515 ;
		RECT	29.13 54.615 29.67 54.825 ;
		RECT	29.13 54.925 29.67 55.02 ;
		RECT	29.13 55.41 29.67 55.51 ;
		RECT	29.13 55.9 29.67 56.005 ;
		RECT	29.13 56.395 29.67 56.485 ;
		RECT	29.13 56.895 29.67 56.985 ;
		RECT	29.13 57.375 29.67 57.48 ;
		RECT	29.13 57.87 29.67 57.97 ;
		RECT	29.13 58.36 29.67 58.465 ;
		RECT	29.13 58.565 29.67 58.755 ;
		RECT	29.13 58.855 29.67 58.955 ;
		RECT	29.13 59.345 29.67 59.445 ;
		RECT	29.13 59.835 29.67 59.94 ;
		RECT	29.13 60.33 29.67 60.43 ;
		RECT	29.13 60.82 29.67 60.925 ;
		RECT	29.13 61.315 29.67 61.415 ;
		RECT	29.13 61.805 29.67 61.905 ;
		RECT	29.13 62.49 29.67 62.7 ;
		RECT	29.13 62.8 29.67 62.89 ;
		RECT	29.13 63.28 29.67 63.375 ;
		RECT	29.13 63.79 29.67 63.86 ;
		RECT	29.13 64.28 29.67 64.35 ;
		RECT	29.13 64.765 29.67 64.825 ;
		RECT	29.13 65.215 29.67 65.35 ;
		RECT	29.13 65.74 29.67 65.81 ;
		RECT	29.13 66.2 29.67 66.35 ;
		RECT	29.13 66.45 29.67 66.64 ;
		RECT	29.13 66.925 29.67 67.115 ;
		RECT	29.13 67.215 29.67 67.32 ;
		RECT	29.13 68.2 29.67 68.305 ;
		RECT	29.13 68.705 29.67 68.915 ;
		RECT	29.67 29.15 30.21 29.34 ;
		RECT	29.67 29.825 30.21 29.925 ;
		RECT	29.67 30.805 30.21 30.91 ;
		RECT	29.67 31.01 30.21 31.2 ;
		RECT	29.67 31.485 30.21 31.675 ;
		RECT	29.67 31.78 30.21 31.93 ;
		RECT	29.67 32.32 30.21 32.385 ;
		RECT	29.67 32.775 30.21 32.88 ;
		RECT	29.67 33.27 30.21 33.37 ;
		RECT	29.67 34.25 30.21 34.355 ;
		RECT	29.67 34.745 30.21 34.845 ;
		RECT	29.67 35.235 30.21 35.34 ;
		RECT	29.67 35.44 30.21 35.63 ;
		RECT	29.67 35.73 30.21 35.83 ;
		RECT	29.67 36.22 30.21 36.325 ;
		RECT	29.67 36.715 30.21 36.815 ;
		RECT	29.67 37.205 30.21 37.305 ;
		RECT	29.67 37.695 30.21 37.8 ;
		RECT	29.67 38.19 30.21 38.29 ;
		RECT	29.67 38.68 30.21 38.78 ;
		RECT	29.67 39.17 30.21 39.275 ;
		RECT	29.67 39.375 30.21 39.565 ;
		RECT	29.67 39.665 30.21 39.765 ;
		RECT	29.67 40.155 30.21 40.26 ;
		RECT	29.67 40.65 30.21 40.75 ;
		RECT	29.67 41.14 30.21 41.23 ;
		RECT	29.67 41.64 30.21 41.735 ;
		RECT	29.67 42.125 30.21 42.225 ;
		RECT	29.67 42.615 30.21 42.72 ;
		RECT	29.67 43.11 30.21 43.2 ;
		RECT	29.67 43.3 30.21 43.51 ;
		RECT	29.67 43.61 30.21 43.705 ;
		RECT	29.67 44.095 30.21 44.2 ;
		RECT	29.67 44.59 30.21 44.685 ;
		RECT	29.67 45.075 30.21 45.18 ;
		RECT	29.67 45.57 30.21 45.655 ;
		RECT	29.67 46.055 30.21 46.265 ;
		RECT	29.67 46.38 30.21 46.57 ;
		RECT	29.67 47.245 30.21 47.435 ;
		RECT	29.67 48.03 30.21 48.13 ;
		RECT	29.67 48.52 30.21 48.62 ;
		RECT	29.67 49.01 30.21 49.115 ;
		RECT	29.67 49.505 30.21 49.605 ;
		RECT	29.67 49.995 30.21 50.1 ;
		RECT	29.67 50.69 30.21 50.88 ;
		RECT	29.67 51.495 30.21 51.685 ;
		RECT	29.67 51.83 30.21 52.04 ;
		RECT	29.67 52.47 30.21 52.555 ;
		RECT	29.67 52.945 30.21 53.05 ;
		RECT	29.67 53.44 30.21 53.545 ;
		RECT	29.67 53.935 30.21 54.025 ;
		RECT	29.67 54.435 30.21 54.515 ;
		RECT	29.67 54.615 30.21 54.825 ;
		RECT	29.67 54.925 30.21 55.02 ;
		RECT	29.67 55.41 30.21 55.51 ;
		RECT	29.67 55.9 30.21 56.005 ;
		RECT	29.67 56.395 30.21 56.485 ;
		RECT	29.67 56.895 30.21 56.985 ;
		RECT	29.67 57.375 30.21 57.48 ;
		RECT	29.67 57.87 30.21 57.97 ;
		RECT	29.67 58.36 30.21 58.465 ;
		RECT	29.67 58.565 30.21 58.755 ;
		RECT	29.67 58.855 30.21 58.955 ;
		RECT	29.67 59.345 30.21 59.445 ;
		RECT	29.67 59.835 30.21 59.94 ;
		RECT	29.67 60.33 30.21 60.43 ;
		RECT	29.67 60.82 30.21 60.925 ;
		RECT	29.67 61.315 30.21 61.415 ;
		RECT	29.67 61.805 30.21 61.905 ;
		RECT	29.67 62.49 30.21 62.7 ;
		RECT	29.67 62.8 30.21 62.89 ;
		RECT	29.67 63.28 30.21 63.375 ;
		RECT	29.67 63.79 30.21 63.86 ;
		RECT	29.67 64.28 30.21 64.35 ;
		RECT	29.67 64.765 30.21 64.825 ;
		RECT	29.67 65.215 30.21 65.35 ;
		RECT	29.67 65.74 30.21 65.81 ;
		RECT	29.67 66.2 30.21 66.35 ;
		RECT	29.67 66.45 30.21 66.64 ;
		RECT	29.67 66.925 30.21 67.115 ;
		RECT	29.67 67.215 30.21 67.32 ;
		RECT	29.67 68.2 30.21 68.305 ;
		RECT	29.67 68.705 30.21 68.915 ;
		RECT	30.21 29.15 30.75 29.34 ;
		RECT	30.21 29.825 30.75 29.925 ;
		RECT	30.21 30.805 30.75 30.91 ;
		RECT	30.21 31.01 30.75 31.2 ;
		RECT	30.21 31.485 30.75 31.675 ;
		RECT	30.21 31.78 30.75 31.93 ;
		RECT	30.21 32.32 30.75 32.385 ;
		RECT	30.21 32.775 30.75 32.88 ;
		RECT	30.21 33.27 30.75 33.37 ;
		RECT	30.21 34.25 30.75 34.355 ;
		RECT	30.21 34.745 30.75 34.845 ;
		RECT	30.21 35.235 30.75 35.34 ;
		RECT	30.21 35.44 30.75 35.63 ;
		RECT	30.21 35.73 30.75 35.83 ;
		RECT	30.21 36.22 30.75 36.325 ;
		RECT	30.21 36.715 30.75 36.815 ;
		RECT	30.21 37.205 30.75 37.305 ;
		RECT	30.21 37.695 30.75 37.8 ;
		RECT	30.21 38.19 30.75 38.29 ;
		RECT	30.21 38.68 30.75 38.78 ;
		RECT	30.21 39.17 30.75 39.275 ;
		RECT	30.21 39.375 30.75 39.565 ;
		RECT	30.21 39.665 30.75 39.765 ;
		RECT	30.21 40.155 30.75 40.26 ;
		RECT	30.21 40.65 30.75 40.75 ;
		RECT	30.21 41.14 30.75 41.23 ;
		RECT	30.21 41.64 30.75 41.735 ;
		RECT	30.21 42.125 30.75 42.225 ;
		RECT	30.21 42.615 30.75 42.72 ;
		RECT	30.21 43.11 30.75 43.2 ;
		RECT	30.21 43.3 30.75 43.51 ;
		RECT	30.21 43.61 30.75 43.705 ;
		RECT	30.21 44.095 30.75 44.2 ;
		RECT	30.21 44.59 30.75 44.685 ;
		RECT	30.21 45.075 30.75 45.18 ;
		RECT	30.21 45.57 30.75 45.655 ;
		RECT	30.21 46.055 30.75 46.265 ;
		RECT	30.21 46.38 30.75 46.57 ;
		RECT	30.21 47.245 30.75 47.435 ;
		RECT	30.21 48.03 30.75 48.13 ;
		RECT	30.21 48.52 30.75 48.62 ;
		RECT	30.21 49.01 30.75 49.115 ;
		RECT	30.21 49.505 30.75 49.605 ;
		RECT	30.21 49.995 30.75 50.1 ;
		RECT	30.21 50.69 30.75 50.88 ;
		RECT	30.21 51.495 30.75 51.685 ;
		RECT	30.21 51.83 30.75 52.04 ;
		RECT	30.21 52.47 30.75 52.555 ;
		RECT	30.21 52.945 30.75 53.05 ;
		RECT	30.21 53.44 30.75 53.545 ;
		RECT	30.21 53.935 30.75 54.025 ;
		RECT	30.21 54.435 30.75 54.515 ;
		RECT	30.21 54.615 30.75 54.825 ;
		RECT	30.21 54.925 30.75 55.02 ;
		RECT	30.21 55.41 30.75 55.51 ;
		RECT	30.21 55.9 30.75 56.005 ;
		RECT	30.21 56.395 30.75 56.485 ;
		RECT	30.21 56.895 30.75 56.985 ;
		RECT	30.21 57.375 30.75 57.48 ;
		RECT	30.21 57.87 30.75 57.97 ;
		RECT	30.21 58.36 30.75 58.465 ;
		RECT	30.21 58.565 30.75 58.755 ;
		RECT	30.21 58.855 30.75 58.955 ;
		RECT	30.21 59.345 30.75 59.445 ;
		RECT	30.21 59.835 30.75 59.94 ;
		RECT	30.21 60.33 30.75 60.43 ;
		RECT	30.21 60.82 30.75 60.925 ;
		RECT	30.21 61.315 30.75 61.415 ;
		RECT	30.21 61.805 30.75 61.905 ;
		RECT	30.21 62.49 30.75 62.7 ;
		RECT	30.21 62.8 30.75 62.89 ;
		RECT	30.21 63.28 30.75 63.375 ;
		RECT	30.21 63.79 30.75 63.86 ;
		RECT	30.21 64.28 30.75 64.35 ;
		RECT	30.21 64.765 30.75 64.825 ;
		RECT	30.21 65.215 30.75 65.35 ;
		RECT	30.21 65.74 30.75 65.81 ;
		RECT	30.21 66.2 30.75 66.35 ;
		RECT	30.21 66.45 30.75 66.64 ;
		RECT	30.21 66.925 30.75 67.115 ;
		RECT	30.21 67.215 30.75 67.32 ;
		RECT	30.21 68.2 30.75 68.305 ;
		RECT	30.21 68.705 30.75 68.915 ;
		RECT	30.75 29.15 31.29 29.34 ;
		RECT	30.75 29.825 31.29 29.925 ;
		RECT	30.75 30.805 31.29 30.91 ;
		RECT	30.75 31.01 31.29 31.2 ;
		RECT	30.75 31.485 31.29 31.675 ;
		RECT	30.75 31.78 31.29 31.93 ;
		RECT	30.75 32.32 31.29 32.385 ;
		RECT	30.75 32.775 31.29 32.88 ;
		RECT	30.75 33.27 31.29 33.37 ;
		RECT	30.75 34.25 31.29 34.355 ;
		RECT	30.75 34.745 31.29 34.845 ;
		RECT	30.75 35.235 31.29 35.34 ;
		RECT	30.75 35.44 31.29 35.63 ;
		RECT	30.75 35.73 31.29 35.83 ;
		RECT	30.75 36.22 31.29 36.325 ;
		RECT	30.75 36.715 31.29 36.815 ;
		RECT	30.75 37.205 31.29 37.305 ;
		RECT	30.75 37.695 31.29 37.8 ;
		RECT	30.75 38.19 31.29 38.29 ;
		RECT	30.75 38.68 31.29 38.78 ;
		RECT	30.75 39.17 31.29 39.275 ;
		RECT	30.75 39.375 31.29 39.565 ;
		RECT	30.75 39.665 31.29 39.765 ;
		RECT	30.75 40.155 31.29 40.26 ;
		RECT	30.75 40.65 31.29 40.75 ;
		RECT	30.75 41.14 31.29 41.23 ;
		RECT	30.75 41.64 31.29 41.735 ;
		RECT	30.75 42.125 31.29 42.225 ;
		RECT	30.75 42.615 31.29 42.72 ;
		RECT	30.75 43.11 31.29 43.2 ;
		RECT	30.75 43.3 31.29 43.51 ;
		RECT	30.75 43.61 31.29 43.705 ;
		RECT	30.75 44.095 31.29 44.2 ;
		RECT	30.75 44.59 31.29 44.685 ;
		RECT	30.75 45.075 31.29 45.18 ;
		RECT	30.75 45.57 31.29 45.655 ;
		RECT	30.75 46.055 31.29 46.265 ;
		RECT	30.75 46.38 31.29 46.57 ;
		RECT	30.75 47.245 31.29 47.435 ;
		RECT	30.75 48.03 31.29 48.13 ;
		RECT	30.75 48.52 31.29 48.62 ;
		RECT	30.75 49.01 31.29 49.115 ;
		RECT	30.75 49.505 31.29 49.605 ;
		RECT	30.75 49.995 31.29 50.1 ;
		RECT	30.75 50.69 31.29 50.88 ;
		RECT	30.75 51.495 31.29 51.685 ;
		RECT	30.75 51.83 31.29 52.04 ;
		RECT	30.75 52.47 31.29 52.555 ;
		RECT	30.75 52.945 31.29 53.05 ;
		RECT	30.75 53.44 31.29 53.545 ;
		RECT	30.75 53.935 31.29 54.025 ;
		RECT	30.75 54.435 31.29 54.515 ;
		RECT	30.75 54.615 31.29 54.825 ;
		RECT	30.75 54.925 31.29 55.02 ;
		RECT	30.75 55.41 31.29 55.51 ;
		RECT	30.75 55.9 31.29 56.005 ;
		RECT	30.75 56.395 31.29 56.485 ;
		RECT	30.75 56.895 31.29 56.985 ;
		RECT	30.75 57.375 31.29 57.48 ;
		RECT	30.75 57.87 31.29 57.97 ;
		RECT	30.75 58.36 31.29 58.465 ;
		RECT	30.75 58.565 31.29 58.755 ;
		RECT	30.75 58.855 31.29 58.955 ;
		RECT	30.75 59.345 31.29 59.445 ;
		RECT	30.75 59.835 31.29 59.94 ;
		RECT	30.75 60.33 31.29 60.43 ;
		RECT	30.75 60.82 31.29 60.925 ;
		RECT	30.75 61.315 31.29 61.415 ;
		RECT	30.75 61.805 31.29 61.905 ;
		RECT	30.75 62.49 31.29 62.7 ;
		RECT	30.75 62.8 31.29 62.89 ;
		RECT	30.75 63.28 31.29 63.375 ;
		RECT	30.75 63.79 31.29 63.86 ;
		RECT	30.75 64.28 31.29 64.35 ;
		RECT	30.75 64.765 31.29 64.825 ;
		RECT	30.75 65.215 31.29 65.35 ;
		RECT	30.75 65.74 31.29 65.81 ;
		RECT	30.75 66.2 31.29 66.35 ;
		RECT	30.75 66.45 31.29 66.64 ;
		RECT	30.75 66.925 31.29 67.115 ;
		RECT	30.75 67.215 31.29 67.32 ;
		RECT	30.75 68.2 31.29 68.305 ;
		RECT	30.75 68.705 31.29 68.915 ;
		RECT	31.29 29.15 31.83 29.34 ;
		RECT	31.29 29.825 31.83 29.925 ;
		RECT	31.29 30.805 31.83 30.91 ;
		RECT	31.29 31.01 31.83 31.2 ;
		RECT	31.29 31.485 31.83 31.675 ;
		RECT	31.29 31.78 31.83 31.93 ;
		RECT	31.29 32.32 31.83 32.385 ;
		RECT	31.29 32.775 31.83 32.88 ;
		RECT	31.29 33.27 31.83 33.37 ;
		RECT	31.29 34.25 31.83 34.355 ;
		RECT	31.29 34.745 31.83 34.845 ;
		RECT	31.29 35.235 31.83 35.34 ;
		RECT	31.29 35.44 31.83 35.63 ;
		RECT	31.29 35.73 31.83 35.83 ;
		RECT	31.29 36.22 31.83 36.325 ;
		RECT	31.29 36.715 31.83 36.815 ;
		RECT	31.29 37.205 31.83 37.305 ;
		RECT	31.29 37.695 31.83 37.8 ;
		RECT	31.29 38.19 31.83 38.29 ;
		RECT	31.29 38.68 31.83 38.78 ;
		RECT	31.29 39.17 31.83 39.275 ;
		RECT	31.29 39.375 31.83 39.565 ;
		RECT	31.29 39.665 31.83 39.765 ;
		RECT	31.29 40.155 31.83 40.26 ;
		RECT	31.29 40.65 31.83 40.75 ;
		RECT	31.29 41.14 31.83 41.23 ;
		RECT	31.29 41.64 31.83 41.735 ;
		RECT	31.29 42.125 31.83 42.225 ;
		RECT	31.29 42.615 31.83 42.72 ;
		RECT	31.29 43.11 31.83 43.2 ;
		RECT	31.29 43.3 31.83 43.51 ;
		RECT	31.29 43.61 31.83 43.705 ;
		RECT	31.29 44.095 31.83 44.2 ;
		RECT	31.29 44.59 31.83 44.685 ;
		RECT	31.29 45.075 31.83 45.18 ;
		RECT	31.29 45.57 31.83 45.655 ;
		RECT	31.29 46.055 31.83 46.265 ;
		RECT	31.29 46.38 31.83 46.57 ;
		RECT	31.29 47.245 31.83 47.435 ;
		RECT	31.29 48.03 31.83 48.13 ;
		RECT	31.29 48.52 31.83 48.62 ;
		RECT	31.29 49.01 31.83 49.115 ;
		RECT	31.29 49.505 31.83 49.605 ;
		RECT	31.29 49.995 31.83 50.1 ;
		RECT	31.29 50.69 31.83 50.88 ;
		RECT	31.29 51.495 31.83 51.685 ;
		RECT	31.29 51.83 31.83 52.04 ;
		RECT	31.29 52.47 31.83 52.555 ;
		RECT	31.29 52.945 31.83 53.05 ;
		RECT	31.29 53.44 31.83 53.545 ;
		RECT	31.29 53.935 31.83 54.025 ;
		RECT	31.29 54.435 31.83 54.515 ;
		RECT	31.29 54.615 31.83 54.825 ;
		RECT	31.29 54.925 31.83 55.02 ;
		RECT	31.29 55.41 31.83 55.51 ;
		RECT	31.29 55.9 31.83 56.005 ;
		RECT	31.29 56.395 31.83 56.485 ;
		RECT	31.29 56.895 31.83 56.985 ;
		RECT	31.29 57.375 31.83 57.48 ;
		RECT	31.29 57.87 31.83 57.97 ;
		RECT	31.29 58.36 31.83 58.465 ;
		RECT	31.29 58.565 31.83 58.755 ;
		RECT	31.29 58.855 31.83 58.955 ;
		RECT	31.29 59.345 31.83 59.445 ;
		RECT	31.29 59.835 31.83 59.94 ;
		RECT	31.29 60.33 31.83 60.43 ;
		RECT	31.29 60.82 31.83 60.925 ;
		RECT	31.29 61.315 31.83 61.415 ;
		RECT	31.29 61.805 31.83 61.905 ;
		RECT	31.29 62.49 31.83 62.7 ;
		RECT	31.29 62.8 31.83 62.89 ;
		RECT	31.29 63.28 31.83 63.375 ;
		RECT	31.29 63.79 31.83 63.86 ;
		RECT	31.29 64.28 31.83 64.35 ;
		RECT	31.29 64.765 31.83 64.825 ;
		RECT	31.29 65.215 31.83 65.35 ;
		RECT	31.29 65.74 31.83 65.81 ;
		RECT	31.29 66.2 31.83 66.35 ;
		RECT	31.29 66.45 31.83 66.64 ;
		RECT	31.29 66.925 31.83 67.115 ;
		RECT	31.29 67.215 31.83 67.32 ;
		RECT	31.29 68.2 31.83 68.305 ;
		RECT	31.29 68.705 31.83 68.915 ;
		RECT	31.83 29.15 32.37 29.34 ;
		RECT	31.83 29.825 32.37 29.925 ;
		RECT	31.83 30.805 32.37 30.91 ;
		RECT	31.83 31.01 32.37 31.2 ;
		RECT	31.83 31.485 32.37 31.675 ;
		RECT	31.83 31.78 32.37 31.93 ;
		RECT	31.83 32.32 32.37 32.385 ;
		RECT	31.83 32.775 32.37 32.88 ;
		RECT	31.83 33.27 32.37 33.37 ;
		RECT	31.83 34.25 32.37 34.355 ;
		RECT	31.83 34.745 32.37 34.845 ;
		RECT	31.83 35.235 32.37 35.34 ;
		RECT	31.83 35.44 32.37 35.63 ;
		RECT	31.83 35.73 32.37 35.83 ;
		RECT	31.83 36.22 32.37 36.325 ;
		RECT	31.83 36.715 32.37 36.815 ;
		RECT	31.83 37.205 32.37 37.305 ;
		RECT	31.83 37.695 32.37 37.8 ;
		RECT	31.83 38.19 32.37 38.29 ;
		RECT	31.83 38.68 32.37 38.78 ;
		RECT	31.83 39.17 32.37 39.275 ;
		RECT	31.83 39.375 32.37 39.565 ;
		RECT	31.83 39.665 32.37 39.765 ;
		RECT	31.83 40.155 32.37 40.26 ;
		RECT	31.83 40.65 32.37 40.75 ;
		RECT	31.83 41.14 32.37 41.23 ;
		RECT	31.83 41.64 32.37 41.735 ;
		RECT	31.83 42.125 32.37 42.225 ;
		RECT	31.83 42.615 32.37 42.72 ;
		RECT	31.83 43.11 32.37 43.2 ;
		RECT	31.83 43.3 32.37 43.51 ;
		RECT	31.83 43.61 32.37 43.705 ;
		RECT	31.83 44.095 32.37 44.2 ;
		RECT	31.83 44.59 32.37 44.685 ;
		RECT	31.83 45.075 32.37 45.18 ;
		RECT	31.83 45.57 32.37 45.655 ;
		RECT	31.83 46.055 32.37 46.265 ;
		RECT	31.83 46.38 32.37 46.57 ;
		RECT	31.83 47.245 32.37 47.435 ;
		RECT	31.83 48.03 32.37 48.13 ;
		RECT	31.83 48.52 32.37 48.62 ;
		RECT	31.83 49.01 32.37 49.115 ;
		RECT	31.83 49.505 32.37 49.605 ;
		RECT	31.83 49.995 32.37 50.1 ;
		RECT	31.83 50.69 32.37 50.88 ;
		RECT	31.83 51.495 32.37 51.685 ;
		RECT	31.83 51.83 32.37 52.04 ;
		RECT	31.83 52.47 32.37 52.555 ;
		RECT	31.83 52.945 32.37 53.05 ;
		RECT	31.83 53.44 32.37 53.545 ;
		RECT	31.83 53.935 32.37 54.025 ;
		RECT	31.83 54.435 32.37 54.515 ;
		RECT	31.83 54.615 32.37 54.825 ;
		RECT	31.83 54.925 32.37 55.02 ;
		RECT	31.83 55.41 32.37 55.51 ;
		RECT	31.83 55.9 32.37 56.005 ;
		RECT	31.83 56.395 32.37 56.485 ;
		RECT	31.83 56.895 32.37 56.985 ;
		RECT	31.83 57.375 32.37 57.48 ;
		RECT	31.83 57.87 32.37 57.97 ;
		RECT	31.83 58.36 32.37 58.465 ;
		RECT	31.83 58.565 32.37 58.755 ;
		RECT	31.83 58.855 32.37 58.955 ;
		RECT	31.83 59.345 32.37 59.445 ;
		RECT	31.83 59.835 32.37 59.94 ;
		RECT	31.83 60.33 32.37 60.43 ;
		RECT	31.83 60.82 32.37 60.925 ;
		RECT	31.83 61.315 32.37 61.415 ;
		RECT	31.83 61.805 32.37 61.905 ;
		RECT	31.83 62.49 32.37 62.7 ;
		RECT	31.83 62.8 32.37 62.89 ;
		RECT	31.83 63.28 32.37 63.375 ;
		RECT	31.83 63.79 32.37 63.86 ;
		RECT	31.83 64.28 32.37 64.35 ;
		RECT	31.83 64.765 32.37 64.825 ;
		RECT	31.83 65.215 32.37 65.35 ;
		RECT	31.83 65.74 32.37 65.81 ;
		RECT	31.83 66.2 32.37 66.35 ;
		RECT	31.83 66.45 32.37 66.64 ;
		RECT	31.83 66.925 32.37 67.115 ;
		RECT	31.83 67.215 32.37 67.32 ;
		RECT	31.83 68.2 32.37 68.305 ;
		RECT	31.83 68.705 32.37 68.915 ;
		RECT	32.37 29.15 32.91 29.34 ;
		RECT	32.37 29.825 32.91 29.925 ;
		RECT	32.37 30.805 32.91 30.91 ;
		RECT	32.37 31.01 32.91 31.2 ;
		RECT	32.37 31.485 32.91 31.675 ;
		RECT	32.37 31.78 32.91 31.93 ;
		RECT	32.37 32.32 32.91 32.385 ;
		RECT	32.37 32.775 32.91 32.88 ;
		RECT	32.37 33.27 32.91 33.37 ;
		RECT	32.37 34.25 32.91 34.355 ;
		RECT	32.37 34.745 32.91 34.845 ;
		RECT	32.37 35.235 32.91 35.34 ;
		RECT	32.37 35.44 32.91 35.63 ;
		RECT	32.37 35.73 32.91 35.83 ;
		RECT	32.37 36.22 32.91 36.325 ;
		RECT	32.37 36.715 32.91 36.815 ;
		RECT	32.37 37.205 32.91 37.305 ;
		RECT	32.37 37.695 32.91 37.8 ;
		RECT	32.37 38.19 32.91 38.29 ;
		RECT	32.37 38.68 32.91 38.78 ;
		RECT	32.37 39.17 32.91 39.275 ;
		RECT	32.37 39.375 32.91 39.565 ;
		RECT	32.37 39.665 32.91 39.765 ;
		RECT	32.37 40.155 32.91 40.26 ;
		RECT	32.37 40.65 32.91 40.75 ;
		RECT	32.37 41.14 32.91 41.23 ;
		RECT	32.37 41.64 32.91 41.735 ;
		RECT	32.37 42.125 32.91 42.225 ;
		RECT	32.37 42.615 32.91 42.72 ;
		RECT	32.37 43.11 32.91 43.2 ;
		RECT	32.37 43.3 32.91 43.51 ;
		RECT	32.37 43.61 32.91 43.705 ;
		RECT	32.37 44.095 32.91 44.2 ;
		RECT	32.37 44.59 32.91 44.685 ;
		RECT	32.37 45.075 32.91 45.18 ;
		RECT	32.37 45.57 32.91 45.655 ;
		RECT	32.37 46.055 32.91 46.265 ;
		RECT	32.37 46.38 32.91 46.57 ;
		RECT	32.37 47.245 32.91 47.435 ;
		RECT	32.37 48.03 32.91 48.13 ;
		RECT	32.37 48.52 32.91 48.62 ;
		RECT	32.37 49.01 32.91 49.115 ;
		RECT	32.37 49.505 32.91 49.605 ;
		RECT	32.37 49.995 32.91 50.1 ;
		RECT	32.37 50.69 32.91 50.88 ;
		RECT	32.37 51.495 32.91 51.685 ;
		RECT	32.37 51.83 32.91 52.04 ;
		RECT	32.37 52.47 32.91 52.555 ;
		RECT	32.37 52.945 32.91 53.05 ;
		RECT	32.37 53.44 32.91 53.545 ;
		RECT	32.37 53.935 32.91 54.025 ;
		RECT	32.37 54.435 32.91 54.515 ;
		RECT	32.37 54.615 32.91 54.825 ;
		RECT	32.37 54.925 32.91 55.02 ;
		RECT	32.37 55.41 32.91 55.51 ;
		RECT	32.37 55.9 32.91 56.005 ;
		RECT	32.37 56.395 32.91 56.485 ;
		RECT	32.37 56.895 32.91 56.985 ;
		RECT	32.37 57.375 32.91 57.48 ;
		RECT	32.37 57.87 32.91 57.97 ;
		RECT	32.37 58.36 32.91 58.465 ;
		RECT	32.37 58.565 32.91 58.755 ;
		RECT	32.37 58.855 32.91 58.955 ;
		RECT	32.37 59.345 32.91 59.445 ;
		RECT	32.37 59.835 32.91 59.94 ;
		RECT	32.37 60.33 32.91 60.43 ;
		RECT	32.37 60.82 32.91 60.925 ;
		RECT	32.37 61.315 32.91 61.415 ;
		RECT	32.37 61.805 32.91 61.905 ;
		RECT	32.37 62.49 32.91 62.7 ;
		RECT	32.37 62.8 32.91 62.89 ;
		RECT	32.37 63.28 32.91 63.375 ;
		RECT	32.37 63.79 32.91 63.86 ;
		RECT	32.37 64.28 32.91 64.35 ;
		RECT	32.37 64.765 32.91 64.825 ;
		RECT	32.37 65.215 32.91 65.35 ;
		RECT	32.37 65.74 32.91 65.81 ;
		RECT	32.37 66.2 32.91 66.35 ;
		RECT	32.37 66.45 32.91 66.64 ;
		RECT	32.37 66.925 32.91 67.115 ;
		RECT	32.37 67.215 32.91 67.32 ;
		RECT	32.37 68.2 32.91 68.305 ;
		RECT	32.37 68.705 32.91 68.915 ;
		RECT	32.91 29.15 33.45 29.34 ;
		RECT	32.91 29.825 33.45 29.925 ;
		RECT	32.91 30.805 33.45 30.91 ;
		RECT	32.91 31.01 33.45 31.2 ;
		RECT	32.91 31.485 33.45 31.675 ;
		RECT	32.91 31.78 33.45 31.93 ;
		RECT	32.91 32.32 33.45 32.385 ;
		RECT	32.91 32.775 33.45 32.88 ;
		RECT	32.91 33.27 33.45 33.37 ;
		RECT	32.91 34.25 33.45 34.355 ;
		RECT	32.91 34.745 33.45 34.845 ;
		RECT	32.91 35.235 33.45 35.34 ;
		RECT	32.91 35.44 33.45 35.63 ;
		RECT	32.91 35.73 33.45 35.83 ;
		RECT	32.91 36.22 33.45 36.325 ;
		RECT	32.91 36.715 33.45 36.815 ;
		RECT	32.91 37.205 33.45 37.305 ;
		RECT	32.91 37.695 33.45 37.8 ;
		RECT	32.91 38.19 33.45 38.29 ;
		RECT	32.91 38.68 33.45 38.78 ;
		RECT	32.91 39.17 33.45 39.275 ;
		RECT	32.91 39.375 33.45 39.565 ;
		RECT	32.91 39.665 33.45 39.765 ;
		RECT	32.91 40.155 33.45 40.26 ;
		RECT	32.91 40.65 33.45 40.75 ;
		RECT	32.91 41.14 33.45 41.23 ;
		RECT	32.91 41.64 33.45 41.735 ;
		RECT	32.91 42.125 33.45 42.225 ;
		RECT	32.91 42.615 33.45 42.72 ;
		RECT	32.91 43.11 33.45 43.2 ;
		RECT	32.91 43.3 33.45 43.51 ;
		RECT	32.91 43.61 33.45 43.705 ;
		RECT	32.91 44.095 33.45 44.2 ;
		RECT	32.91 44.59 33.45 44.685 ;
		RECT	32.91 45.075 33.45 45.18 ;
		RECT	32.91 45.57 33.45 45.655 ;
		RECT	32.91 46.055 33.45 46.265 ;
		RECT	32.91 46.38 33.45 46.57 ;
		RECT	32.91 47.245 33.45 47.435 ;
		RECT	32.91 48.03 33.45 48.13 ;
		RECT	32.91 48.52 33.45 48.62 ;
		RECT	32.91 49.01 33.45 49.115 ;
		RECT	32.91 49.505 33.45 49.605 ;
		RECT	32.91 49.995 33.45 50.1 ;
		RECT	32.91 50.69 33.45 50.88 ;
		RECT	32.91 51.495 33.45 51.685 ;
		RECT	32.91 51.83 33.45 52.04 ;
		RECT	32.91 52.47 33.45 52.555 ;
		RECT	32.91 52.945 33.45 53.05 ;
		RECT	32.91 53.44 33.45 53.545 ;
		RECT	32.91 53.935 33.45 54.025 ;
		RECT	32.91 54.435 33.45 54.515 ;
		RECT	32.91 54.615 33.45 54.825 ;
		RECT	32.91 54.925 33.45 55.02 ;
		RECT	32.91 55.41 33.45 55.51 ;
		RECT	32.91 55.9 33.45 56.005 ;
		RECT	32.91 56.395 33.45 56.485 ;
		RECT	32.91 56.895 33.45 56.985 ;
		RECT	32.91 57.375 33.45 57.48 ;
		RECT	32.91 57.87 33.45 57.97 ;
		RECT	32.91 58.36 33.45 58.465 ;
		RECT	32.91 58.565 33.45 58.755 ;
		RECT	32.91 58.855 33.45 58.955 ;
		RECT	32.91 59.345 33.45 59.445 ;
		RECT	32.91 59.835 33.45 59.94 ;
		RECT	32.91 60.33 33.45 60.43 ;
		RECT	32.91 60.82 33.45 60.925 ;
		RECT	32.91 61.315 33.45 61.415 ;
		RECT	32.91 61.805 33.45 61.905 ;
		RECT	32.91 62.49 33.45 62.7 ;
		RECT	32.91 62.8 33.45 62.89 ;
		RECT	32.91 63.28 33.45 63.375 ;
		RECT	32.91 63.79 33.45 63.86 ;
		RECT	32.91 64.28 33.45 64.35 ;
		RECT	32.91 64.765 33.45 64.825 ;
		RECT	32.91 65.215 33.45 65.35 ;
		RECT	32.91 65.74 33.45 65.81 ;
		RECT	32.91 66.2 33.45 66.35 ;
		RECT	32.91 66.45 33.45 66.64 ;
		RECT	32.91 66.925 33.45 67.115 ;
		RECT	32.91 67.215 33.45 67.32 ;
		RECT	32.91 68.2 33.45 68.305 ;
		RECT	32.91 68.705 33.45 68.915 ;
		RECT	33.45 29.15 33.99 29.34 ;
		RECT	33.45 29.825 33.99 29.925 ;
		RECT	33.45 30.805 33.99 30.91 ;
		RECT	33.45 31.01 33.99 31.2 ;
		RECT	33.45 31.485 33.99 31.675 ;
		RECT	33.45 31.78 33.99 31.93 ;
		RECT	33.45 32.32 33.99 32.385 ;
		RECT	33.45 32.775 33.99 32.88 ;
		RECT	33.45 33.27 33.99 33.37 ;
		RECT	33.45 34.25 33.99 34.355 ;
		RECT	33.45 34.745 33.99 34.845 ;
		RECT	33.45 35.235 33.99 35.34 ;
		RECT	33.45 35.44 33.99 35.63 ;
		RECT	33.45 35.73 33.99 35.83 ;
		RECT	33.45 36.22 33.99 36.325 ;
		RECT	33.45 36.715 33.99 36.815 ;
		RECT	33.45 37.205 33.99 37.305 ;
		RECT	33.45 37.695 33.99 37.8 ;
		RECT	33.45 38.19 33.99 38.29 ;
		RECT	33.45 38.68 33.99 38.78 ;
		RECT	33.45 39.17 33.99 39.275 ;
		RECT	33.45 39.375 33.99 39.565 ;
		RECT	33.45 39.665 33.99 39.765 ;
		RECT	33.45 40.155 33.99 40.26 ;
		RECT	33.45 40.65 33.99 40.75 ;
		RECT	33.45 41.14 33.99 41.23 ;
		RECT	33.45 41.64 33.99 41.735 ;
		RECT	33.45 42.125 33.99 42.225 ;
		RECT	33.45 42.615 33.99 42.72 ;
		RECT	33.45 43.11 33.99 43.2 ;
		RECT	33.45 43.3 33.99 43.51 ;
		RECT	33.45 43.61 33.99 43.705 ;
		RECT	33.45 44.095 33.99 44.2 ;
		RECT	33.45 44.59 33.99 44.685 ;
		RECT	33.45 45.075 33.99 45.18 ;
		RECT	33.45 45.57 33.99 45.655 ;
		RECT	33.45 46.055 33.99 46.265 ;
		RECT	33.45 46.38 33.99 46.57 ;
		RECT	33.45 47.245 33.99 47.435 ;
		RECT	33.45 48.03 33.99 48.13 ;
		RECT	33.45 48.52 33.99 48.62 ;
		RECT	33.45 49.01 33.99 49.115 ;
		RECT	33.45 49.505 33.99 49.605 ;
		RECT	33.45 49.995 33.99 50.1 ;
		RECT	33.45 50.69 33.99 50.88 ;
		RECT	33.45 51.495 33.99 51.685 ;
		RECT	33.45 51.83 33.99 52.04 ;
		RECT	33.45 52.47 33.99 52.555 ;
		RECT	33.45 52.945 33.99 53.05 ;
		RECT	33.45 53.44 33.99 53.545 ;
		RECT	33.45 53.935 33.99 54.025 ;
		RECT	33.45 54.435 33.99 54.515 ;
		RECT	33.45 54.615 33.99 54.825 ;
		RECT	33.45 54.925 33.99 55.02 ;
		RECT	33.45 55.41 33.99 55.51 ;
		RECT	33.45 55.9 33.99 56.005 ;
		RECT	33.45 56.395 33.99 56.485 ;
		RECT	33.45 56.895 33.99 56.985 ;
		RECT	33.45 57.375 33.99 57.48 ;
		RECT	33.45 57.87 33.99 57.97 ;
		RECT	33.45 58.36 33.99 58.465 ;
		RECT	33.45 58.565 33.99 58.755 ;
		RECT	33.45 58.855 33.99 58.955 ;
		RECT	33.45 59.345 33.99 59.445 ;
		RECT	33.45 59.835 33.99 59.94 ;
		RECT	33.45 60.33 33.99 60.43 ;
		RECT	33.45 60.82 33.99 60.925 ;
		RECT	33.45 61.315 33.99 61.415 ;
		RECT	33.45 61.805 33.99 61.905 ;
		RECT	33.45 62.49 33.99 62.7 ;
		RECT	33.45 62.8 33.99 62.89 ;
		RECT	33.45 63.28 33.99 63.375 ;
		RECT	33.45 63.79 33.99 63.86 ;
		RECT	33.45 64.28 33.99 64.35 ;
		RECT	33.45 64.765 33.99 64.825 ;
		RECT	33.45 65.215 33.99 65.35 ;
		RECT	33.45 65.74 33.99 65.81 ;
		RECT	33.45 66.2 33.99 66.35 ;
		RECT	33.45 66.45 33.99 66.64 ;
		RECT	33.45 66.925 33.99 67.115 ;
		RECT	33.45 67.215 33.99 67.32 ;
		RECT	33.45 68.2 33.99 68.305 ;
		RECT	33.45 68.705 33.99 68.915 ;
		RECT	33.99 29.15 34.53 29.34 ;
		RECT	33.99 29.825 34.53 29.925 ;
		RECT	33.99 30.805 34.53 30.91 ;
		RECT	33.99 31.01 34.53 31.2 ;
		RECT	33.99 31.485 34.53 31.675 ;
		RECT	33.99 31.78 34.53 31.93 ;
		RECT	33.99 32.32 34.53 32.385 ;
		RECT	33.99 32.775 34.53 32.88 ;
		RECT	33.99 33.27 34.53 33.37 ;
		RECT	33.99 34.25 34.53 34.355 ;
		RECT	33.99 34.745 34.53 34.845 ;
		RECT	33.99 35.235 34.53 35.34 ;
		RECT	33.99 35.44 34.53 35.63 ;
		RECT	33.99 35.73 34.53 35.83 ;
		RECT	33.99 36.22 34.53 36.325 ;
		RECT	33.99 36.715 34.53 36.815 ;
		RECT	33.99 37.205 34.53 37.305 ;
		RECT	33.99 37.695 34.53 37.8 ;
		RECT	33.99 38.19 34.53 38.29 ;
		RECT	33.99 38.68 34.53 38.78 ;
		RECT	33.99 39.17 34.53 39.275 ;
		RECT	33.99 39.375 34.53 39.565 ;
		RECT	33.99 39.665 34.53 39.765 ;
		RECT	33.99 40.155 34.53 40.26 ;
		RECT	33.99 40.65 34.53 40.75 ;
		RECT	33.99 41.14 34.53 41.23 ;
		RECT	33.99 41.64 34.53 41.735 ;
		RECT	33.99 42.125 34.53 42.225 ;
		RECT	33.99 42.615 34.53 42.72 ;
		RECT	33.99 43.11 34.53 43.2 ;
		RECT	33.99 43.3 34.53 43.51 ;
		RECT	33.99 43.61 34.53 43.705 ;
		RECT	33.99 44.095 34.53 44.2 ;
		RECT	33.99 44.59 34.53 44.685 ;
		RECT	33.99 45.075 34.53 45.18 ;
		RECT	33.99 45.57 34.53 45.655 ;
		RECT	33.99 46.055 34.53 46.265 ;
		RECT	33.99 46.38 34.53 46.57 ;
		RECT	33.99 47.245 34.53 47.435 ;
		RECT	33.99 48.03 34.53 48.13 ;
		RECT	33.99 48.52 34.53 48.62 ;
		RECT	33.99 49.01 34.53 49.115 ;
		RECT	33.99 49.505 34.53 49.605 ;
		RECT	33.99 49.995 34.53 50.1 ;
		RECT	33.99 50.69 34.53 50.88 ;
		RECT	33.99 51.495 34.53 51.685 ;
		RECT	33.99 51.83 34.53 52.04 ;
		RECT	33.99 52.47 34.53 52.555 ;
		RECT	33.99 52.945 34.53 53.05 ;
		RECT	33.99 53.44 34.53 53.545 ;
		RECT	33.99 53.935 34.53 54.025 ;
		RECT	33.99 54.435 34.53 54.515 ;
		RECT	33.99 54.615 34.53 54.825 ;
		RECT	33.99 54.925 34.53 55.02 ;
		RECT	33.99 55.41 34.53 55.51 ;
		RECT	33.99 55.9 34.53 56.005 ;
		RECT	33.99 56.395 34.53 56.485 ;
		RECT	33.99 56.895 34.53 56.985 ;
		RECT	33.99 57.375 34.53 57.48 ;
		RECT	33.99 57.87 34.53 57.97 ;
		RECT	33.99 58.36 34.53 58.465 ;
		RECT	33.99 58.565 34.53 58.755 ;
		RECT	33.99 58.855 34.53 58.955 ;
		RECT	33.99 59.345 34.53 59.445 ;
		RECT	33.99 59.835 34.53 59.94 ;
		RECT	33.99 60.33 34.53 60.43 ;
		RECT	33.99 60.82 34.53 60.925 ;
		RECT	33.99 61.315 34.53 61.415 ;
		RECT	33.99 61.805 34.53 61.905 ;
		RECT	33.99 62.49 34.53 62.7 ;
		RECT	33.99 62.8 34.53 62.89 ;
		RECT	33.99 63.28 34.53 63.375 ;
		RECT	33.99 63.79 34.53 63.86 ;
		RECT	33.99 64.28 34.53 64.35 ;
		RECT	33.99 64.765 34.53 64.825 ;
		RECT	33.99 65.215 34.53 65.35 ;
		RECT	33.99 65.74 34.53 65.81 ;
		RECT	33.99 66.2 34.53 66.35 ;
		RECT	33.99 66.45 34.53 66.64 ;
		RECT	33.99 66.925 34.53 67.115 ;
		RECT	33.99 67.215 34.53 67.32 ;
		RECT	33.99 68.2 34.53 68.305 ;
		RECT	33.99 68.705 34.53 68.915 ;
		RECT	34.53 29.15 35.07 29.34 ;
		RECT	34.53 29.825 35.07 29.925 ;
		RECT	34.53 30.805 35.07 30.91 ;
		RECT	34.53 31.01 35.07 31.2 ;
		RECT	34.53 31.485 35.07 31.675 ;
		RECT	34.53 31.78 35.07 31.93 ;
		RECT	34.53 32.32 35.07 32.385 ;
		RECT	34.53 32.775 35.07 32.88 ;
		RECT	34.53 33.27 35.07 33.37 ;
		RECT	34.53 34.25 35.07 34.355 ;
		RECT	34.53 34.745 35.07 34.845 ;
		RECT	34.53 35.235 35.07 35.34 ;
		RECT	34.53 35.44 35.07 35.63 ;
		RECT	34.53 35.73 35.07 35.83 ;
		RECT	34.53 36.22 35.07 36.325 ;
		RECT	34.53 36.715 35.07 36.815 ;
		RECT	34.53 37.205 35.07 37.305 ;
		RECT	34.53 37.695 35.07 37.8 ;
		RECT	34.53 38.19 35.07 38.29 ;
		RECT	34.53 38.68 35.07 38.78 ;
		RECT	34.53 39.17 35.07 39.275 ;
		RECT	34.53 39.375 35.07 39.565 ;
		RECT	34.53 39.665 35.07 39.765 ;
		RECT	34.53 40.155 35.07 40.26 ;
		RECT	34.53 40.65 35.07 40.75 ;
		RECT	34.53 41.14 35.07 41.23 ;
		RECT	34.53 41.64 35.07 41.735 ;
		RECT	34.53 42.125 35.07 42.225 ;
		RECT	34.53 42.615 35.07 42.72 ;
		RECT	34.53 43.11 35.07 43.2 ;
		RECT	34.53 43.3 35.07 43.51 ;
		RECT	34.53 43.61 35.07 43.705 ;
		RECT	34.53 44.095 35.07 44.2 ;
		RECT	34.53 44.59 35.07 44.685 ;
		RECT	34.53 45.075 35.07 45.18 ;
		RECT	34.53 45.57 35.07 45.655 ;
		RECT	34.53 46.055 35.07 46.265 ;
		RECT	34.53 46.38 35.07 46.57 ;
		RECT	34.53 47.245 35.07 47.435 ;
		RECT	34.53 48.03 35.07 48.13 ;
		RECT	34.53 48.52 35.07 48.62 ;
		RECT	34.53 49.01 35.07 49.115 ;
		RECT	34.53 49.505 35.07 49.605 ;
		RECT	34.53 49.995 35.07 50.1 ;
		RECT	34.53 50.69 35.07 50.88 ;
		RECT	34.53 51.495 35.07 51.685 ;
		RECT	34.53 51.83 35.07 52.04 ;
		RECT	34.53 52.47 35.07 52.555 ;
		RECT	34.53 52.945 35.07 53.05 ;
		RECT	34.53 53.44 35.07 53.545 ;
		RECT	34.53 53.935 35.07 54.025 ;
		RECT	34.53 54.435 35.07 54.515 ;
		RECT	34.53 54.615 35.07 54.825 ;
		RECT	34.53 54.925 35.07 55.02 ;
		RECT	34.53 55.41 35.07 55.51 ;
		RECT	34.53 55.9 35.07 56.005 ;
		RECT	34.53 56.395 35.07 56.485 ;
		RECT	34.53 56.895 35.07 56.985 ;
		RECT	34.53 57.375 35.07 57.48 ;
		RECT	34.53 57.87 35.07 57.97 ;
		RECT	34.53 58.36 35.07 58.465 ;
		RECT	34.53 58.565 35.07 58.755 ;
		RECT	34.53 58.855 35.07 58.955 ;
		RECT	34.53 59.345 35.07 59.445 ;
		RECT	34.53 59.835 35.07 59.94 ;
		RECT	34.53 60.33 35.07 60.43 ;
		RECT	34.53 60.82 35.07 60.925 ;
		RECT	34.53 61.315 35.07 61.415 ;
		RECT	34.53 61.805 35.07 61.905 ;
		RECT	34.53 62.49 35.07 62.7 ;
		RECT	34.53 62.8 35.07 62.89 ;
		RECT	34.53 63.28 35.07 63.375 ;
		RECT	34.53 63.79 35.07 63.86 ;
		RECT	34.53 64.28 35.07 64.35 ;
		RECT	34.53 64.765 35.07 64.825 ;
		RECT	34.53 65.215 35.07 65.35 ;
		RECT	34.53 65.74 35.07 65.81 ;
		RECT	34.53 66.2 35.07 66.35 ;
		RECT	34.53 66.45 35.07 66.64 ;
		RECT	34.53 66.925 35.07 67.115 ;
		RECT	34.53 67.215 35.07 67.32 ;
		RECT	34.53 68.2 35.07 68.305 ;
		RECT	34.53 68.705 35.07 68.915 ;
		RECT	35.07 29.15 35.61 29.34 ;
		RECT	35.07 29.825 35.61 29.925 ;
		RECT	35.07 30.805 35.61 30.91 ;
		RECT	35.07 31.01 35.61 31.2 ;
		RECT	35.07 31.485 35.61 31.675 ;
		RECT	35.07 31.78 35.61 31.93 ;
		RECT	35.07 32.32 35.61 32.385 ;
		RECT	35.07 32.775 35.61 32.88 ;
		RECT	35.07 33.27 35.61 33.37 ;
		RECT	35.07 34.25 35.61 34.355 ;
		RECT	35.07 34.745 35.61 34.845 ;
		RECT	35.07 35.235 35.61 35.34 ;
		RECT	35.07 35.44 35.61 35.63 ;
		RECT	35.07 35.73 35.61 35.83 ;
		RECT	35.07 36.22 35.61 36.325 ;
		RECT	35.07 36.715 35.61 36.815 ;
		RECT	35.07 37.205 35.61 37.305 ;
		RECT	35.07 37.695 35.61 37.8 ;
		RECT	35.07 38.19 35.61 38.29 ;
		RECT	35.07 38.68 35.61 38.78 ;
		RECT	35.07 39.17 35.61 39.275 ;
		RECT	35.07 39.375 35.61 39.565 ;
		RECT	35.07 39.665 35.61 39.765 ;
		RECT	35.07 40.155 35.61 40.26 ;
		RECT	35.07 40.65 35.61 40.75 ;
		RECT	35.07 41.14 35.61 41.23 ;
		RECT	35.07 41.64 35.61 41.735 ;
		RECT	35.07 42.125 35.61 42.225 ;
		RECT	35.07 42.615 35.61 42.72 ;
		RECT	35.07 43.11 35.61 43.2 ;
		RECT	35.07 43.3 35.61 43.51 ;
		RECT	35.07 43.61 35.61 43.705 ;
		RECT	35.07 44.095 35.61 44.2 ;
		RECT	35.07 44.59 35.61 44.685 ;
		RECT	35.07 45.075 35.61 45.18 ;
		RECT	35.07 45.57 35.61 45.655 ;
		RECT	35.07 46.055 35.61 46.265 ;
		RECT	35.07 46.38 35.61 46.57 ;
		RECT	35.07 47.245 35.61 47.435 ;
		RECT	35.07 48.03 35.61 48.13 ;
		RECT	35.07 48.52 35.61 48.62 ;
		RECT	35.07 49.01 35.61 49.115 ;
		RECT	35.07 49.505 35.61 49.605 ;
		RECT	35.07 49.995 35.61 50.1 ;
		RECT	35.07 50.69 35.61 50.88 ;
		RECT	35.07 51.495 35.61 51.685 ;
		RECT	35.07 51.83 35.61 52.04 ;
		RECT	35.07 52.47 35.61 52.555 ;
		RECT	35.07 52.945 35.61 53.05 ;
		RECT	35.07 53.44 35.61 53.545 ;
		RECT	35.07 53.935 35.61 54.025 ;
		RECT	35.07 54.435 35.61 54.515 ;
		RECT	35.07 54.615 35.61 54.825 ;
		RECT	35.07 54.925 35.61 55.02 ;
		RECT	35.07 55.41 35.61 55.51 ;
		RECT	35.07 55.9 35.61 56.005 ;
		RECT	35.07 56.395 35.61 56.485 ;
		RECT	35.07 56.895 35.61 56.985 ;
		RECT	35.07 57.375 35.61 57.48 ;
		RECT	35.07 57.87 35.61 57.97 ;
		RECT	35.07 58.36 35.61 58.465 ;
		RECT	35.07 58.565 35.61 58.755 ;
		RECT	35.07 58.855 35.61 58.955 ;
		RECT	35.07 59.345 35.61 59.445 ;
		RECT	35.07 59.835 35.61 59.94 ;
		RECT	35.07 60.33 35.61 60.43 ;
		RECT	35.07 60.82 35.61 60.925 ;
		RECT	35.07 61.315 35.61 61.415 ;
		RECT	35.07 61.805 35.61 61.905 ;
		RECT	35.07 62.49 35.61 62.7 ;
		RECT	35.07 62.8 35.61 62.89 ;
		RECT	35.07 63.28 35.61 63.375 ;
		RECT	35.07 63.79 35.61 63.86 ;
		RECT	35.07 64.28 35.61 64.35 ;
		RECT	35.07 64.765 35.61 64.825 ;
		RECT	35.07 65.215 35.61 65.35 ;
		RECT	35.07 65.74 35.61 65.81 ;
		RECT	35.07 66.2 35.61 66.35 ;
		RECT	35.07 66.45 35.61 66.64 ;
		RECT	35.07 66.925 35.61 67.115 ;
		RECT	35.07 67.215 35.61 67.32 ;
		RECT	35.07 68.2 35.61 68.305 ;
		RECT	35.07 68.705 35.61 68.915 ;
		RECT	35.61 29.15 36.15 29.34 ;
		RECT	35.61 29.825 36.15 29.925 ;
		RECT	35.61 30.805 36.15 30.91 ;
		RECT	35.61 31.01 36.15 31.2 ;
		RECT	35.61 31.485 36.15 31.675 ;
		RECT	35.61 31.78 36.15 31.93 ;
		RECT	35.61 32.32 36.15 32.385 ;
		RECT	35.61 32.775 36.15 32.88 ;
		RECT	35.61 33.27 36.15 33.37 ;
		RECT	35.61 34.25 36.15 34.355 ;
		RECT	35.61 34.745 36.15 34.845 ;
		RECT	35.61 35.235 36.15 35.34 ;
		RECT	35.61 35.44 36.15 35.63 ;
		RECT	35.61 35.73 36.15 35.83 ;
		RECT	35.61 36.22 36.15 36.325 ;
		RECT	35.61 36.715 36.15 36.815 ;
		RECT	35.61 37.205 36.15 37.305 ;
		RECT	35.61 37.695 36.15 37.8 ;
		RECT	35.61 38.19 36.15 38.29 ;
		RECT	35.61 38.68 36.15 38.78 ;
		RECT	35.61 39.17 36.15 39.275 ;
		RECT	35.61 39.375 36.15 39.565 ;
		RECT	35.61 39.665 36.15 39.765 ;
		RECT	35.61 40.155 36.15 40.26 ;
		RECT	35.61 40.65 36.15 40.75 ;
		RECT	35.61 41.14 36.15 41.23 ;
		RECT	35.61 41.64 36.15 41.735 ;
		RECT	35.61 42.125 36.15 42.225 ;
		RECT	35.61 42.615 36.15 42.72 ;
		RECT	35.61 43.11 36.15 43.2 ;
		RECT	35.61 43.3 36.15 43.51 ;
		RECT	35.61 43.61 36.15 43.705 ;
		RECT	35.61 44.095 36.15 44.2 ;
		RECT	35.61 44.59 36.15 44.685 ;
		RECT	35.61 45.075 36.15 45.18 ;
		RECT	35.61 45.57 36.15 45.655 ;
		RECT	35.61 46.055 36.15 46.265 ;
		RECT	35.61 46.38 36.15 46.57 ;
		RECT	35.61 47.245 36.15 47.435 ;
		RECT	35.61 48.03 36.15 48.13 ;
		RECT	35.61 48.52 36.15 48.62 ;
		RECT	35.61 49.01 36.15 49.115 ;
		RECT	35.61 49.505 36.15 49.605 ;
		RECT	35.61 49.995 36.15 50.1 ;
		RECT	35.61 50.69 36.15 50.88 ;
		RECT	35.61 51.495 36.15 51.685 ;
		RECT	35.61 51.83 36.15 52.04 ;
		RECT	35.61 52.47 36.15 52.555 ;
		RECT	35.61 52.945 36.15 53.05 ;
		RECT	35.61 53.44 36.15 53.545 ;
		RECT	35.61 53.935 36.15 54.025 ;
		RECT	35.61 54.435 36.15 54.515 ;
		RECT	35.61 54.615 36.15 54.825 ;
		RECT	35.61 54.925 36.15 55.02 ;
		RECT	35.61 55.41 36.15 55.51 ;
		RECT	35.61 55.9 36.15 56.005 ;
		RECT	35.61 56.395 36.15 56.485 ;
		RECT	35.61 56.895 36.15 56.985 ;
		RECT	35.61 57.375 36.15 57.48 ;
		RECT	35.61 57.87 36.15 57.97 ;
		RECT	35.61 58.36 36.15 58.465 ;
		RECT	35.61 58.565 36.15 58.755 ;
		RECT	35.61 58.855 36.15 58.955 ;
		RECT	35.61 59.345 36.15 59.445 ;
		RECT	35.61 59.835 36.15 59.94 ;
		RECT	35.61 60.33 36.15 60.43 ;
		RECT	35.61 60.82 36.15 60.925 ;
		RECT	35.61 61.315 36.15 61.415 ;
		RECT	35.61 61.805 36.15 61.905 ;
		RECT	35.61 62.49 36.15 62.7 ;
		RECT	35.61 62.8 36.15 62.89 ;
		RECT	35.61 63.28 36.15 63.375 ;
		RECT	35.61 63.79 36.15 63.86 ;
		RECT	35.61 64.28 36.15 64.35 ;
		RECT	35.61 64.765 36.15 64.825 ;
		RECT	35.61 65.215 36.15 65.35 ;
		RECT	35.61 65.74 36.15 65.81 ;
		RECT	35.61 66.2 36.15 66.35 ;
		RECT	35.61 66.45 36.15 66.64 ;
		RECT	35.61 66.925 36.15 67.115 ;
		RECT	35.61 67.215 36.15 67.32 ;
		RECT	35.61 68.2 36.15 68.305 ;
		RECT	35.61 68.705 36.15 68.915 ;
		RECT	36.15 29.15 36.69 29.34 ;
		RECT	36.15 29.825 36.69 29.925 ;
		RECT	36.15 30.805 36.69 30.91 ;
		RECT	36.15 31.01 36.69 31.2 ;
		RECT	36.15 31.485 36.69 31.675 ;
		RECT	36.15 31.78 36.69 31.93 ;
		RECT	36.15 32.32 36.69 32.385 ;
		RECT	36.15 32.775 36.69 32.88 ;
		RECT	36.15 33.27 36.69 33.37 ;
		RECT	36.15 34.25 36.69 34.355 ;
		RECT	36.15 34.745 36.69 34.845 ;
		RECT	36.15 35.235 36.69 35.34 ;
		RECT	36.15 35.44 36.69 35.63 ;
		RECT	36.15 35.73 36.69 35.83 ;
		RECT	36.15 36.22 36.69 36.325 ;
		RECT	36.15 36.715 36.69 36.815 ;
		RECT	36.15 37.205 36.69 37.305 ;
		RECT	36.15 37.695 36.69 37.8 ;
		RECT	36.15 38.19 36.69 38.29 ;
		RECT	36.15 38.68 36.69 38.78 ;
		RECT	36.15 39.17 36.69 39.275 ;
		RECT	36.15 39.375 36.69 39.565 ;
		RECT	36.15 39.665 36.69 39.765 ;
		RECT	36.15 40.155 36.69 40.26 ;
		RECT	36.15 40.65 36.69 40.75 ;
		RECT	36.15 41.14 36.69 41.23 ;
		RECT	36.15 41.64 36.69 41.735 ;
		RECT	36.15 42.125 36.69 42.225 ;
		RECT	36.15 42.615 36.69 42.72 ;
		RECT	36.15 43.11 36.69 43.2 ;
		RECT	36.15 43.3 36.69 43.51 ;
		RECT	36.15 43.61 36.69 43.705 ;
		RECT	36.15 44.095 36.69 44.2 ;
		RECT	36.15 44.59 36.69 44.685 ;
		RECT	36.15 45.075 36.69 45.18 ;
		RECT	36.15 45.57 36.69 45.655 ;
		RECT	36.15 46.055 36.69 46.265 ;
		RECT	36.15 46.38 36.69 46.57 ;
		RECT	36.15 47.245 36.69 47.435 ;
		RECT	36.15 48.03 36.69 48.13 ;
		RECT	36.15 48.52 36.69 48.62 ;
		RECT	36.15 49.01 36.69 49.115 ;
		RECT	36.15 49.505 36.69 49.605 ;
		RECT	36.15 49.995 36.69 50.1 ;
		RECT	36.15 50.69 36.69 50.88 ;
		RECT	36.15 51.495 36.69 51.685 ;
		RECT	36.15 51.83 36.69 52.04 ;
		RECT	36.15 52.47 36.69 52.555 ;
		RECT	36.15 52.945 36.69 53.05 ;
		RECT	36.15 53.44 36.69 53.545 ;
		RECT	36.15 53.935 36.69 54.025 ;
		RECT	36.15 54.435 36.69 54.515 ;
		RECT	36.15 54.615 36.69 54.825 ;
		RECT	36.15 54.925 36.69 55.02 ;
		RECT	36.15 55.41 36.69 55.51 ;
		RECT	36.15 55.9 36.69 56.005 ;
		RECT	36.15 56.395 36.69 56.485 ;
		RECT	36.15 56.895 36.69 56.985 ;
		RECT	36.15 57.375 36.69 57.48 ;
		RECT	36.15 57.87 36.69 57.97 ;
		RECT	36.15 58.36 36.69 58.465 ;
		RECT	36.15 58.565 36.69 58.755 ;
		RECT	36.15 58.855 36.69 58.955 ;
		RECT	36.15 59.345 36.69 59.445 ;
		RECT	36.15 59.835 36.69 59.94 ;
		RECT	36.15 60.33 36.69 60.43 ;
		RECT	36.15 60.82 36.69 60.925 ;
		RECT	36.15 61.315 36.69 61.415 ;
		RECT	36.15 61.805 36.69 61.905 ;
		RECT	36.15 62.49 36.69 62.7 ;
		RECT	36.15 62.8 36.69 62.89 ;
		RECT	36.15 63.28 36.69 63.375 ;
		RECT	36.15 63.79 36.69 63.86 ;
		RECT	36.15 64.28 36.69 64.35 ;
		RECT	36.15 64.765 36.69 64.825 ;
		RECT	36.15 65.215 36.69 65.35 ;
		RECT	36.15 65.74 36.69 65.81 ;
		RECT	36.15 66.2 36.69 66.35 ;
		RECT	36.15 66.45 36.69 66.64 ;
		RECT	36.15 66.925 36.69 67.115 ;
		RECT	36.15 67.215 36.69 67.32 ;
		RECT	36.15 68.2 36.69 68.305 ;
		RECT	36.15 68.705 36.69 68.915 ;
		RECT	36.69 29.15 37.23 29.34 ;
		RECT	36.69 29.825 37.23 29.925 ;
		RECT	36.69 30.805 37.23 30.91 ;
		RECT	36.69 31.01 37.23 31.2 ;
		RECT	36.69 31.485 37.23 31.675 ;
		RECT	36.69 31.78 37.23 31.93 ;
		RECT	36.69 32.32 37.23 32.385 ;
		RECT	36.69 32.775 37.23 32.88 ;
		RECT	36.69 33.27 37.23 33.37 ;
		RECT	36.69 34.25 37.23 34.355 ;
		RECT	36.69 34.745 37.23 34.845 ;
		RECT	36.69 35.235 37.23 35.34 ;
		RECT	36.69 35.44 37.23 35.63 ;
		RECT	36.69 35.73 37.23 35.83 ;
		RECT	36.69 36.22 37.23 36.325 ;
		RECT	36.69 36.715 37.23 36.815 ;
		RECT	36.69 37.205 37.23 37.305 ;
		RECT	36.69 37.695 37.23 37.8 ;
		RECT	36.69 38.19 37.23 38.29 ;
		RECT	36.69 38.68 37.23 38.78 ;
		RECT	36.69 39.17 37.23 39.275 ;
		RECT	36.69 39.375 37.23 39.565 ;
		RECT	36.69 39.665 37.23 39.765 ;
		RECT	36.69 40.155 37.23 40.26 ;
		RECT	36.69 40.65 37.23 40.75 ;
		RECT	36.69 41.14 37.23 41.23 ;
		RECT	36.69 41.64 37.23 41.735 ;
		RECT	36.69 42.125 37.23 42.225 ;
		RECT	36.69 42.615 37.23 42.72 ;
		RECT	36.69 43.11 37.23 43.2 ;
		RECT	36.69 43.3 37.23 43.51 ;
		RECT	36.69 43.61 37.23 43.705 ;
		RECT	36.69 44.095 37.23 44.2 ;
		RECT	36.69 44.59 37.23 44.685 ;
		RECT	36.69 45.075 37.23 45.18 ;
		RECT	36.69 45.57 37.23 45.655 ;
		RECT	36.69 46.055 37.23 46.265 ;
		RECT	36.69 46.38 37.23 46.57 ;
		RECT	36.69 47.245 37.23 47.435 ;
		RECT	36.69 48.03 37.23 48.13 ;
		RECT	36.69 48.52 37.23 48.62 ;
		RECT	36.69 49.01 37.23 49.115 ;
		RECT	36.69 49.505 37.23 49.605 ;
		RECT	36.69 49.995 37.23 50.1 ;
		RECT	36.69 50.69 37.23 50.88 ;
		RECT	36.69 51.495 37.23 51.685 ;
		RECT	36.69 51.83 37.23 52.04 ;
		RECT	36.69 52.47 37.23 52.555 ;
		RECT	36.69 52.945 37.23 53.05 ;
		RECT	36.69 53.44 37.23 53.545 ;
		RECT	36.69 53.935 37.23 54.025 ;
		RECT	36.69 54.435 37.23 54.515 ;
		RECT	36.69 54.615 37.23 54.825 ;
		RECT	36.69 54.925 37.23 55.02 ;
		RECT	36.69 55.41 37.23 55.51 ;
		RECT	36.69 55.9 37.23 56.005 ;
		RECT	36.69 56.395 37.23 56.485 ;
		RECT	36.69 56.895 37.23 56.985 ;
		RECT	36.69 57.375 37.23 57.48 ;
		RECT	36.69 57.87 37.23 57.97 ;
		RECT	36.69 58.36 37.23 58.465 ;
		RECT	36.69 58.565 37.23 58.755 ;
		RECT	36.69 58.855 37.23 58.955 ;
		RECT	36.69 59.345 37.23 59.445 ;
		RECT	36.69 59.835 37.23 59.94 ;
		RECT	36.69 60.33 37.23 60.43 ;
		RECT	36.69 60.82 37.23 60.925 ;
		RECT	36.69 61.315 37.23 61.415 ;
		RECT	36.69 61.805 37.23 61.905 ;
		RECT	36.69 62.49 37.23 62.7 ;
		RECT	36.69 62.8 37.23 62.89 ;
		RECT	36.69 63.28 37.23 63.375 ;
		RECT	36.69 63.79 37.23 63.86 ;
		RECT	36.69 64.28 37.23 64.35 ;
		RECT	36.69 64.765 37.23 64.825 ;
		RECT	36.69 65.215 37.23 65.35 ;
		RECT	36.69 65.74 37.23 65.81 ;
		RECT	36.69 66.2 37.23 66.35 ;
		RECT	36.69 66.45 37.23 66.64 ;
		RECT	36.69 66.925 37.23 67.115 ;
		RECT	36.69 67.215 37.23 67.32 ;
		RECT	36.69 68.2 37.23 68.305 ;
		RECT	36.69 68.705 37.23 68.915 ;
		RECT	37.23 29.15 37.77 29.34 ;
		RECT	37.23 29.825 37.77 29.925 ;
		RECT	37.23 30.805 37.77 30.91 ;
		RECT	37.23 31.01 37.77 31.2 ;
		RECT	37.23 31.485 37.77 31.675 ;
		RECT	37.23 31.78 37.77 31.93 ;
		RECT	37.23 32.32 37.77 32.385 ;
		RECT	37.23 32.775 37.77 32.88 ;
		RECT	37.23 33.27 37.77 33.37 ;
		RECT	37.23 34.25 37.77 34.355 ;
		RECT	37.23 34.745 37.77 34.845 ;
		RECT	37.23 35.235 37.77 35.34 ;
		RECT	37.23 35.44 37.77 35.63 ;
		RECT	37.23 35.73 37.77 35.83 ;
		RECT	37.23 36.22 37.77 36.325 ;
		RECT	37.23 36.715 37.77 36.815 ;
		RECT	37.23 37.205 37.77 37.305 ;
		RECT	37.23 37.695 37.77 37.8 ;
		RECT	37.23 38.19 37.77 38.29 ;
		RECT	37.23 38.68 37.77 38.78 ;
		RECT	37.23 39.17 37.77 39.275 ;
		RECT	37.23 39.375 37.77 39.565 ;
		RECT	37.23 39.665 37.77 39.765 ;
		RECT	37.23 40.155 37.77 40.26 ;
		RECT	37.23 40.65 37.77 40.75 ;
		RECT	37.23 41.14 37.77 41.23 ;
		RECT	37.23 41.64 37.77 41.735 ;
		RECT	37.23 42.125 37.77 42.225 ;
		RECT	37.23 42.615 37.77 42.72 ;
		RECT	37.23 43.11 37.77 43.2 ;
		RECT	37.23 43.3 37.77 43.51 ;
		RECT	37.23 43.61 37.77 43.705 ;
		RECT	37.23 44.095 37.77 44.2 ;
		RECT	37.23 44.59 37.77 44.685 ;
		RECT	37.23 45.075 37.77 45.18 ;
		RECT	37.23 45.57 37.77 45.655 ;
		RECT	37.23 46.055 37.77 46.265 ;
		RECT	37.23 46.38 37.77 46.57 ;
		RECT	37.23 47.245 37.77 47.435 ;
		RECT	37.23 48.03 37.77 48.13 ;
		RECT	37.23 48.52 37.77 48.62 ;
		RECT	37.23 49.01 37.77 49.115 ;
		RECT	37.23 49.505 37.77 49.605 ;
		RECT	37.23 49.995 37.77 50.1 ;
		RECT	37.23 50.69 37.77 50.88 ;
		RECT	37.23 51.495 37.77 51.685 ;
		RECT	37.23 51.83 37.77 52.04 ;
		RECT	37.23 52.47 37.77 52.555 ;
		RECT	37.23 52.945 37.77 53.05 ;
		RECT	37.23 53.44 37.77 53.545 ;
		RECT	37.23 53.935 37.77 54.025 ;
		RECT	37.23 54.435 37.77 54.515 ;
		RECT	37.23 54.615 37.77 54.825 ;
		RECT	37.23 54.925 37.77 55.02 ;
		RECT	37.23 55.41 37.77 55.51 ;
		RECT	37.23 55.9 37.77 56.005 ;
		RECT	37.23 56.395 37.77 56.485 ;
		RECT	37.23 56.895 37.77 56.985 ;
		RECT	37.23 57.375 37.77 57.48 ;
		RECT	37.23 57.87 37.77 57.97 ;
		RECT	37.23 58.36 37.77 58.465 ;
		RECT	37.23 58.565 37.77 58.755 ;
		RECT	37.23 58.855 37.77 58.955 ;
		RECT	37.23 59.345 37.77 59.445 ;
		RECT	37.23 59.835 37.77 59.94 ;
		RECT	37.23 60.33 37.77 60.43 ;
		RECT	37.23 60.82 37.77 60.925 ;
		RECT	37.23 61.315 37.77 61.415 ;
		RECT	37.23 61.805 37.77 61.905 ;
		RECT	37.23 62.49 37.77 62.7 ;
		RECT	37.23 62.8 37.77 62.89 ;
		RECT	37.23 63.28 37.77 63.375 ;
		RECT	37.23 63.79 37.77 63.86 ;
		RECT	37.23 64.28 37.77 64.35 ;
		RECT	37.23 64.765 37.77 64.825 ;
		RECT	37.23 65.215 37.77 65.35 ;
		RECT	37.23 65.74 37.77 65.81 ;
		RECT	37.23 66.2 37.77 66.35 ;
		RECT	37.23 66.45 37.77 66.64 ;
		RECT	37.23 66.925 37.77 67.115 ;
		RECT	37.23 67.215 37.77 67.32 ;
		RECT	37.23 68.2 37.77 68.305 ;
		RECT	37.23 68.705 37.77 68.915 ;
		RECT	37.77 29.15 38.31 29.34 ;
		RECT	37.77 29.825 38.31 29.925 ;
		RECT	37.77 30.805 38.31 30.91 ;
		RECT	37.77 31.01 38.31 31.2 ;
		RECT	37.77 31.485 38.31 31.675 ;
		RECT	37.77 31.78 38.31 31.93 ;
		RECT	37.77 32.32 38.31 32.385 ;
		RECT	37.77 32.775 38.31 32.88 ;
		RECT	37.77 33.27 38.31 33.37 ;
		RECT	37.77 34.25 38.31 34.355 ;
		RECT	37.77 34.745 38.31 34.845 ;
		RECT	37.77 35.235 38.31 35.34 ;
		RECT	37.77 35.44 38.31 35.63 ;
		RECT	37.77 35.73 38.31 35.83 ;
		RECT	37.77 36.22 38.31 36.325 ;
		RECT	37.77 36.715 38.31 36.815 ;
		RECT	37.77 37.205 38.31 37.305 ;
		RECT	37.77 37.695 38.31 37.8 ;
		RECT	37.77 38.19 38.31 38.29 ;
		RECT	37.77 38.68 38.31 38.78 ;
		RECT	37.77 39.17 38.31 39.275 ;
		RECT	37.77 39.375 38.31 39.565 ;
		RECT	37.77 39.665 38.31 39.765 ;
		RECT	37.77 40.155 38.31 40.26 ;
		RECT	37.77 40.65 38.31 40.75 ;
		RECT	37.77 41.14 38.31 41.23 ;
		RECT	37.77 41.64 38.31 41.735 ;
		RECT	37.77 42.125 38.31 42.225 ;
		RECT	37.77 42.615 38.31 42.72 ;
		RECT	37.77 43.11 38.31 43.2 ;
		RECT	37.77 43.3 38.31 43.51 ;
		RECT	37.77 43.61 38.31 43.705 ;
		RECT	37.77 44.095 38.31 44.2 ;
		RECT	37.77 44.59 38.31 44.685 ;
		RECT	37.77 45.075 38.31 45.18 ;
		RECT	37.77 45.57 38.31 45.655 ;
		RECT	37.77 46.055 38.31 46.265 ;
		RECT	37.77 46.38 38.31 46.57 ;
		RECT	37.77 47.245 38.31 47.435 ;
		RECT	37.77 48.03 38.31 48.13 ;
		RECT	37.77 48.52 38.31 48.62 ;
		RECT	37.77 49.01 38.31 49.115 ;
		RECT	37.77 49.505 38.31 49.605 ;
		RECT	37.77 49.995 38.31 50.1 ;
		RECT	37.77 50.69 38.31 50.88 ;
		RECT	37.77 51.495 38.31 51.685 ;
		RECT	37.77 51.83 38.31 52.04 ;
		RECT	37.77 52.47 38.31 52.555 ;
		RECT	37.77 52.945 38.31 53.05 ;
		RECT	37.77 53.44 38.31 53.545 ;
		RECT	37.77 53.935 38.31 54.025 ;
		RECT	37.77 54.435 38.31 54.515 ;
		RECT	37.77 54.615 38.31 54.825 ;
		RECT	37.77 54.925 38.31 55.02 ;
		RECT	37.77 55.41 38.31 55.51 ;
		RECT	37.77 55.9 38.31 56.005 ;
		RECT	37.77 56.395 38.31 56.485 ;
		RECT	37.77 56.895 38.31 56.985 ;
		RECT	37.77 57.375 38.31 57.48 ;
		RECT	37.77 57.87 38.31 57.97 ;
		RECT	37.77 58.36 38.31 58.465 ;
		RECT	37.77 58.565 38.31 58.755 ;
		RECT	37.77 58.855 38.31 58.955 ;
		RECT	37.77 59.345 38.31 59.445 ;
		RECT	37.77 59.835 38.31 59.94 ;
		RECT	37.77 60.33 38.31 60.43 ;
		RECT	37.77 60.82 38.31 60.925 ;
		RECT	37.77 61.315 38.31 61.415 ;
		RECT	37.77 61.805 38.31 61.905 ;
		RECT	37.77 62.49 38.31 62.7 ;
		RECT	37.77 62.8 38.31 62.89 ;
		RECT	37.77 63.28 38.31 63.375 ;
		RECT	37.77 63.79 38.31 63.86 ;
		RECT	37.77 64.28 38.31 64.35 ;
		RECT	37.77 64.765 38.31 64.825 ;
		RECT	37.77 65.215 38.31 65.35 ;
		RECT	37.77 65.74 38.31 65.81 ;
		RECT	37.77 66.2 38.31 66.35 ;
		RECT	37.77 66.45 38.31 66.64 ;
		RECT	37.77 66.925 38.31 67.115 ;
		RECT	37.77 67.215 38.31 67.32 ;
		RECT	37.77 68.2 38.31 68.305 ;
		RECT	37.77 68.705 38.31 68.915 ;
		RECT	38.31 29.15 38.85 29.34 ;
		RECT	38.31 29.825 38.85 29.925 ;
		RECT	38.31 30.805 38.85 30.91 ;
		RECT	38.31 31.01 38.85 31.2 ;
		RECT	38.31 31.485 38.85 31.675 ;
		RECT	38.31 31.78 38.85 31.93 ;
		RECT	38.31 32.32 38.85 32.385 ;
		RECT	38.31 32.775 38.85 32.88 ;
		RECT	38.31 33.27 38.85 33.37 ;
		RECT	38.31 34.25 38.85 34.355 ;
		RECT	38.31 34.745 38.85 34.845 ;
		RECT	38.31 35.235 38.85 35.34 ;
		RECT	38.31 35.44 38.85 35.63 ;
		RECT	38.31 35.73 38.85 35.83 ;
		RECT	38.31 36.22 38.85 36.325 ;
		RECT	38.31 36.715 38.85 36.815 ;
		RECT	38.31 37.205 38.85 37.305 ;
		RECT	38.31 37.695 38.85 37.8 ;
		RECT	38.31 38.19 38.85 38.29 ;
		RECT	38.31 38.68 38.85 38.78 ;
		RECT	38.31 39.17 38.85 39.275 ;
		RECT	38.31 39.375 38.85 39.565 ;
		RECT	38.31 39.665 38.85 39.765 ;
		RECT	38.31 40.155 38.85 40.26 ;
		RECT	38.31 40.65 38.85 40.75 ;
		RECT	38.31 41.14 38.85 41.23 ;
		RECT	38.31 41.64 38.85 41.735 ;
		RECT	38.31 42.125 38.85 42.225 ;
		RECT	38.31 42.615 38.85 42.72 ;
		RECT	38.31 43.11 38.85 43.2 ;
		RECT	38.31 43.3 38.85 43.51 ;
		RECT	38.31 43.61 38.85 43.705 ;
		RECT	38.31 44.095 38.85 44.2 ;
		RECT	38.31 44.59 38.85 44.685 ;
		RECT	38.31 45.075 38.85 45.18 ;
		RECT	38.31 45.57 38.85 45.655 ;
		RECT	38.31 46.055 38.85 46.265 ;
		RECT	38.31 46.38 38.85 46.57 ;
		RECT	38.31 47.245 38.85 47.435 ;
		RECT	38.31 48.03 38.85 48.13 ;
		RECT	38.31 48.52 38.85 48.62 ;
		RECT	38.31 49.01 38.85 49.115 ;
		RECT	38.31 49.505 38.85 49.605 ;
		RECT	38.31 49.995 38.85 50.1 ;
		RECT	38.31 50.69 38.85 50.88 ;
		RECT	38.31 51.495 38.85 51.685 ;
		RECT	38.31 51.83 38.85 52.04 ;
		RECT	38.31 52.47 38.85 52.555 ;
		RECT	38.31 52.945 38.85 53.05 ;
		RECT	38.31 53.44 38.85 53.545 ;
		RECT	38.31 53.935 38.85 54.025 ;
		RECT	38.31 54.435 38.85 54.515 ;
		RECT	38.31 54.615 38.85 54.825 ;
		RECT	38.31 54.925 38.85 55.02 ;
		RECT	38.31 55.41 38.85 55.51 ;
		RECT	38.31 55.9 38.85 56.005 ;
		RECT	38.31 56.395 38.85 56.485 ;
		RECT	38.31 56.895 38.85 56.985 ;
		RECT	38.31 57.375 38.85 57.48 ;
		RECT	38.31 57.87 38.85 57.97 ;
		RECT	38.31 58.36 38.85 58.465 ;
		RECT	38.31 58.565 38.85 58.755 ;
		RECT	38.31 58.855 38.85 58.955 ;
		RECT	38.31 59.345 38.85 59.445 ;
		RECT	38.31 59.835 38.85 59.94 ;
		RECT	38.31 60.33 38.85 60.43 ;
		RECT	38.31 60.82 38.85 60.925 ;
		RECT	38.31 61.315 38.85 61.415 ;
		RECT	38.31 61.805 38.85 61.905 ;
		RECT	38.31 62.49 38.85 62.7 ;
		RECT	38.31 62.8 38.85 62.89 ;
		RECT	38.31 63.28 38.85 63.375 ;
		RECT	38.31 63.79 38.85 63.86 ;
		RECT	38.31 64.28 38.85 64.35 ;
		RECT	38.31 64.765 38.85 64.825 ;
		RECT	38.31 65.215 38.85 65.35 ;
		RECT	38.31 65.74 38.85 65.81 ;
		RECT	38.31 66.2 38.85 66.35 ;
		RECT	38.31 66.45 38.85 66.64 ;
		RECT	38.31 66.925 38.85 67.115 ;
		RECT	38.31 67.215 38.85 67.32 ;
		RECT	38.31 68.2 38.85 68.305 ;
		RECT	38.31 68.705 38.85 68.915 ;
		RECT	38.85 29.15 39.39 29.34 ;
		RECT	38.85 29.825 39.39 29.925 ;
		RECT	38.85 30.805 39.39 30.91 ;
		RECT	38.85 31.01 39.39 31.2 ;
		RECT	38.85 31.485 39.39 31.675 ;
		RECT	38.85 31.78 39.39 31.93 ;
		RECT	38.85 32.32 39.39 32.385 ;
		RECT	38.85 32.775 39.39 32.88 ;
		RECT	38.85 33.27 39.39 33.37 ;
		RECT	38.85 34.25 39.39 34.355 ;
		RECT	38.85 34.745 39.39 34.845 ;
		RECT	38.85 35.235 39.39 35.34 ;
		RECT	38.85 35.44 39.39 35.63 ;
		RECT	38.85 35.73 39.39 35.83 ;
		RECT	38.85 36.22 39.39 36.325 ;
		RECT	38.85 36.715 39.39 36.815 ;
		RECT	38.85 37.205 39.39 37.305 ;
		RECT	38.85 37.695 39.39 37.8 ;
		RECT	38.85 38.19 39.39 38.29 ;
		RECT	38.85 38.68 39.39 38.78 ;
		RECT	38.85 39.17 39.39 39.275 ;
		RECT	38.85 39.375 39.39 39.565 ;
		RECT	38.85 39.665 39.39 39.765 ;
		RECT	38.85 40.155 39.39 40.26 ;
		RECT	38.85 40.65 39.39 40.75 ;
		RECT	38.85 41.14 39.39 41.23 ;
		RECT	38.85 41.64 39.39 41.735 ;
		RECT	38.85 42.125 39.39 42.225 ;
		RECT	38.85 42.615 39.39 42.72 ;
		RECT	38.85 43.11 39.39 43.2 ;
		RECT	38.85 43.3 39.39 43.51 ;
		RECT	38.85 43.61 39.39 43.705 ;
		RECT	38.85 44.095 39.39 44.2 ;
		RECT	38.85 44.59 39.39 44.685 ;
		RECT	38.85 45.075 39.39 45.18 ;
		RECT	38.85 45.57 39.39 45.655 ;
		RECT	38.85 46.055 39.39 46.265 ;
		RECT	38.85 46.38 39.39 46.57 ;
		RECT	38.85 47.245 39.39 47.435 ;
		RECT	38.85 48.03 39.39 48.13 ;
		RECT	38.85 48.52 39.39 48.62 ;
		RECT	38.85 49.01 39.39 49.115 ;
		RECT	38.85 49.505 39.39 49.605 ;
		RECT	38.85 49.995 39.39 50.1 ;
		RECT	38.85 50.69 39.39 50.88 ;
		RECT	38.85 51.495 39.39 51.685 ;
		RECT	38.85 51.83 39.39 52.04 ;
		RECT	38.85 52.47 39.39 52.555 ;
		RECT	38.85 52.945 39.39 53.05 ;
		RECT	38.85 53.44 39.39 53.545 ;
		RECT	38.85 53.935 39.39 54.025 ;
		RECT	38.85 54.435 39.39 54.515 ;
		RECT	38.85 54.615 39.39 54.825 ;
		RECT	38.85 54.925 39.39 55.02 ;
		RECT	38.85 55.41 39.39 55.51 ;
		RECT	38.85 55.9 39.39 56.005 ;
		RECT	38.85 56.395 39.39 56.485 ;
		RECT	38.85 56.895 39.39 56.985 ;
		RECT	38.85 57.375 39.39 57.48 ;
		RECT	38.85 57.87 39.39 57.97 ;
		RECT	38.85 58.36 39.39 58.465 ;
		RECT	38.85 58.565 39.39 58.755 ;
		RECT	38.85 58.855 39.39 58.955 ;
		RECT	38.85 59.345 39.39 59.445 ;
		RECT	38.85 59.835 39.39 59.94 ;
		RECT	38.85 60.33 39.39 60.43 ;
		RECT	38.85 60.82 39.39 60.925 ;
		RECT	38.85 61.315 39.39 61.415 ;
		RECT	38.85 61.805 39.39 61.905 ;
		RECT	38.85 62.49 39.39 62.7 ;
		RECT	38.85 62.8 39.39 62.89 ;
		RECT	38.85 63.28 39.39 63.375 ;
		RECT	38.85 63.79 39.39 63.86 ;
		RECT	38.85 64.28 39.39 64.35 ;
		RECT	38.85 64.765 39.39 64.825 ;
		RECT	38.85 65.215 39.39 65.35 ;
		RECT	38.85 65.74 39.39 65.81 ;
		RECT	38.85 66.2 39.39 66.35 ;
		RECT	38.85 66.45 39.39 66.64 ;
		RECT	38.85 66.925 39.39 67.115 ;
		RECT	38.85 67.215 39.39 67.32 ;
		RECT	38.85 68.2 39.39 68.305 ;
		RECT	38.85 68.705 39.39 68.915 ;
		RECT	39.39 29.15 39.93 29.34 ;
		RECT	39.39 29.825 39.93 29.925 ;
		RECT	39.39 30.805 39.93 30.91 ;
		RECT	39.39 31.01 39.93 31.2 ;
		RECT	39.39 31.485 39.93 31.675 ;
		RECT	39.39 31.78 39.93 31.93 ;
		RECT	39.39 32.32 39.93 32.385 ;
		RECT	39.39 32.775 39.93 32.88 ;
		RECT	39.39 33.27 39.93 33.37 ;
		RECT	39.39 34.25 39.93 34.355 ;
		RECT	39.39 34.745 39.93 34.845 ;
		RECT	39.39 35.235 39.93 35.34 ;
		RECT	39.39 35.44 39.93 35.63 ;
		RECT	39.39 35.73 39.93 35.83 ;
		RECT	39.39 36.22 39.93 36.325 ;
		RECT	39.39 36.715 39.93 36.815 ;
		RECT	39.39 37.205 39.93 37.305 ;
		RECT	39.39 37.695 39.93 37.8 ;
		RECT	39.39 38.19 39.93 38.29 ;
		RECT	39.39 38.68 39.93 38.78 ;
		RECT	39.39 39.17 39.93 39.275 ;
		RECT	39.39 39.375 39.93 39.565 ;
		RECT	39.39 39.665 39.93 39.765 ;
		RECT	39.39 40.155 39.93 40.26 ;
		RECT	39.39 40.65 39.93 40.75 ;
		RECT	39.39 41.14 39.93 41.23 ;
		RECT	39.39 41.64 39.93 41.735 ;
		RECT	39.39 42.125 39.93 42.225 ;
		RECT	39.39 42.615 39.93 42.72 ;
		RECT	39.39 43.11 39.93 43.2 ;
		RECT	39.39 43.3 39.93 43.51 ;
		RECT	39.39 43.61 39.93 43.705 ;
		RECT	39.39 44.095 39.93 44.2 ;
		RECT	39.39 44.59 39.93 44.685 ;
		RECT	39.39 45.075 39.93 45.18 ;
		RECT	39.39 45.57 39.93 45.655 ;
		RECT	39.39 46.055 39.93 46.265 ;
		RECT	39.39 46.38 39.93 46.57 ;
		RECT	39.39 47.245 39.93 47.435 ;
		RECT	39.39 48.03 39.93 48.13 ;
		RECT	39.39 48.52 39.93 48.62 ;
		RECT	39.39 49.01 39.93 49.115 ;
		RECT	39.39 49.505 39.93 49.605 ;
		RECT	39.39 49.995 39.93 50.1 ;
		RECT	39.39 50.69 39.93 50.88 ;
		RECT	39.39 51.495 39.93 51.685 ;
		RECT	39.39 51.83 39.93 52.04 ;
		RECT	39.39 52.47 39.93 52.555 ;
		RECT	39.39 52.945 39.93 53.05 ;
		RECT	39.39 53.44 39.93 53.545 ;
		RECT	39.39 53.935 39.93 54.025 ;
		RECT	39.39 54.435 39.93 54.515 ;
		RECT	39.39 54.615 39.93 54.825 ;
		RECT	39.39 54.925 39.93 55.02 ;
		RECT	39.39 55.41 39.93 55.51 ;
		RECT	39.39 55.9 39.93 56.005 ;
		RECT	39.39 56.395 39.93 56.485 ;
		RECT	39.39 56.895 39.93 56.985 ;
		RECT	39.39 57.375 39.93 57.48 ;
		RECT	39.39 57.87 39.93 57.97 ;
		RECT	39.39 58.36 39.93 58.465 ;
		RECT	39.39 58.565 39.93 58.755 ;
		RECT	39.39 58.855 39.93 58.955 ;
		RECT	39.39 59.345 39.93 59.445 ;
		RECT	39.39 59.835 39.93 59.94 ;
		RECT	39.39 60.33 39.93 60.43 ;
		RECT	39.39 60.82 39.93 60.925 ;
		RECT	39.39 61.315 39.93 61.415 ;
		RECT	39.39 61.805 39.93 61.905 ;
		RECT	39.39 62.49 39.93 62.7 ;
		RECT	39.39 62.8 39.93 62.89 ;
		RECT	39.39 63.28 39.93 63.375 ;
		RECT	39.39 63.79 39.93 63.86 ;
		RECT	39.39 64.28 39.93 64.35 ;
		RECT	39.39 64.765 39.93 64.825 ;
		RECT	39.39 65.215 39.93 65.35 ;
		RECT	39.39 65.74 39.93 65.81 ;
		RECT	39.39 66.2 39.93 66.35 ;
		RECT	39.39 66.45 39.93 66.64 ;
		RECT	39.39 66.925 39.93 67.115 ;
		RECT	39.39 67.215 39.93 67.32 ;
		RECT	39.39 68.2 39.93 68.305 ;
		RECT	39.39 68.705 39.93 68.915 ;
		RECT	39.93 29.15 40.47 29.34 ;
		RECT	39.93 29.825 40.47 29.925 ;
		RECT	39.93 30.805 40.47 30.91 ;
		RECT	39.93 31.01 40.47 31.2 ;
		RECT	39.93 31.485 40.47 31.675 ;
		RECT	39.93 31.78 40.47 31.93 ;
		RECT	39.93 32.32 40.47 32.385 ;
		RECT	39.93 32.775 40.47 32.88 ;
		RECT	39.93 33.27 40.47 33.37 ;
		RECT	39.93 34.25 40.47 34.355 ;
		RECT	39.93 34.745 40.47 34.845 ;
		RECT	39.93 35.235 40.47 35.34 ;
		RECT	39.93 35.44 40.47 35.63 ;
		RECT	39.93 35.73 40.47 35.83 ;
		RECT	39.93 36.22 40.47 36.325 ;
		RECT	39.93 36.715 40.47 36.815 ;
		RECT	39.93 37.205 40.47 37.305 ;
		RECT	39.93 37.695 40.47 37.8 ;
		RECT	39.93 38.19 40.47 38.29 ;
		RECT	39.93 38.68 40.47 38.78 ;
		RECT	39.93 39.17 40.47 39.275 ;
		RECT	39.93 39.375 40.47 39.565 ;
		RECT	39.93 39.665 40.47 39.765 ;
		RECT	39.93 40.155 40.47 40.26 ;
		RECT	39.93 40.65 40.47 40.75 ;
		RECT	39.93 41.14 40.47 41.23 ;
		RECT	39.93 41.64 40.47 41.735 ;
		RECT	39.93 42.125 40.47 42.225 ;
		RECT	39.93 42.615 40.47 42.72 ;
		RECT	39.93 43.11 40.47 43.2 ;
		RECT	39.93 43.3 40.47 43.51 ;
		RECT	39.93 43.61 40.47 43.705 ;
		RECT	39.93 44.095 40.47 44.2 ;
		RECT	39.93 44.59 40.47 44.685 ;
		RECT	39.93 45.075 40.47 45.18 ;
		RECT	39.93 45.57 40.47 45.655 ;
		RECT	39.93 46.055 40.47 46.265 ;
		RECT	39.93 46.38 40.47 46.57 ;
		RECT	39.93 47.245 40.47 47.435 ;
		RECT	39.93 48.03 40.47 48.13 ;
		RECT	39.93 48.52 40.47 48.62 ;
		RECT	39.93 49.01 40.47 49.115 ;
		RECT	39.93 49.505 40.47 49.605 ;
		RECT	39.93 49.995 40.47 50.1 ;
		RECT	39.93 50.69 40.47 50.88 ;
		RECT	39.93 51.495 40.47 51.685 ;
		RECT	39.93 51.83 40.47 52.04 ;
		RECT	39.93 52.47 40.47 52.555 ;
		RECT	39.93 52.945 40.47 53.05 ;
		RECT	39.93 53.44 40.47 53.545 ;
		RECT	39.93 53.935 40.47 54.025 ;
		RECT	39.93 54.435 40.47 54.515 ;
		RECT	39.93 54.615 40.47 54.825 ;
		RECT	39.93 54.925 40.47 55.02 ;
		RECT	39.93 55.41 40.47 55.51 ;
		RECT	39.93 55.9 40.47 56.005 ;
		RECT	39.93 56.395 40.47 56.485 ;
		RECT	39.93 56.895 40.47 56.985 ;
		RECT	39.93 57.375 40.47 57.48 ;
		RECT	39.93 57.87 40.47 57.97 ;
		RECT	39.93 58.36 40.47 58.465 ;
		RECT	39.93 58.565 40.47 58.755 ;
		RECT	39.93 58.855 40.47 58.955 ;
		RECT	39.93 59.345 40.47 59.445 ;
		RECT	39.93 59.835 40.47 59.94 ;
		RECT	39.93 60.33 40.47 60.43 ;
		RECT	39.93 60.82 40.47 60.925 ;
		RECT	39.93 61.315 40.47 61.415 ;
		RECT	39.93 61.805 40.47 61.905 ;
		RECT	39.93 62.49 40.47 62.7 ;
		RECT	39.93 62.8 40.47 62.89 ;
		RECT	39.93 63.28 40.47 63.375 ;
		RECT	39.93 63.79 40.47 63.86 ;
		RECT	39.93 64.28 40.47 64.35 ;
		RECT	39.93 64.765 40.47 64.825 ;
		RECT	39.93 65.215 40.47 65.35 ;
		RECT	39.93 65.74 40.47 65.81 ;
		RECT	39.93 66.2 40.47 66.35 ;
		RECT	39.93 66.45 40.47 66.64 ;
		RECT	39.93 66.925 40.47 67.115 ;
		RECT	39.93 67.215 40.47 67.32 ;
		RECT	39.93 68.2 40.47 68.305 ;
		RECT	39.93 68.705 40.47 68.915 ;
		RECT	40.47 29.15 41.01 29.34 ;
		RECT	40.47 29.825 41.01 29.925 ;
		RECT	40.47 30.805 41.01 30.91 ;
		RECT	40.47 31.01 41.01 31.2 ;
		RECT	40.47 31.485 41.01 31.675 ;
		RECT	40.47 31.78 41.01 31.93 ;
		RECT	40.47 32.32 41.01 32.385 ;
		RECT	40.47 32.775 41.01 32.88 ;
		RECT	40.47 33.27 41.01 33.37 ;
		RECT	40.47 34.25 41.01 34.355 ;
		RECT	40.47 34.745 41.01 34.845 ;
		RECT	40.47 35.235 41.01 35.34 ;
		RECT	40.47 35.44 41.01 35.63 ;
		RECT	40.47 35.73 41.01 35.83 ;
		RECT	40.47 36.22 41.01 36.325 ;
		RECT	40.47 36.715 41.01 36.815 ;
		RECT	40.47 37.205 41.01 37.305 ;
		RECT	40.47 37.695 41.01 37.8 ;
		RECT	40.47 38.19 41.01 38.29 ;
		RECT	40.47 38.68 41.01 38.78 ;
		RECT	40.47 39.17 41.01 39.275 ;
		RECT	40.47 39.375 41.01 39.565 ;
		RECT	40.47 39.665 41.01 39.765 ;
		RECT	40.47 40.155 41.01 40.26 ;
		RECT	40.47 40.65 41.01 40.75 ;
		RECT	40.47 41.14 41.01 41.23 ;
		RECT	40.47 41.64 41.01 41.735 ;
		RECT	40.47 42.125 41.01 42.225 ;
		RECT	40.47 42.615 41.01 42.72 ;
		RECT	40.47 43.11 41.01 43.2 ;
		RECT	40.47 43.3 41.01 43.51 ;
		RECT	40.47 43.61 41.01 43.705 ;
		RECT	40.47 44.095 41.01 44.2 ;
		RECT	40.47 44.59 41.01 44.685 ;
		RECT	40.47 45.075 41.01 45.18 ;
		RECT	40.47 45.57 41.01 45.655 ;
		RECT	40.47 46.055 41.01 46.265 ;
		RECT	40.47 46.38 41.01 46.57 ;
		RECT	40.47 47.245 41.01 47.435 ;
		RECT	40.47 48.03 41.01 48.13 ;
		RECT	40.47 48.52 41.01 48.62 ;
		RECT	40.47 49.01 41.01 49.115 ;
		RECT	40.47 49.505 41.01 49.605 ;
		RECT	40.47 49.995 41.01 50.1 ;
		RECT	40.47 50.69 41.01 50.88 ;
		RECT	40.47 51.495 41.01 51.685 ;
		RECT	40.47 51.83 41.01 52.04 ;
		RECT	40.47 52.47 41.01 52.555 ;
		RECT	40.47 52.945 41.01 53.05 ;
		RECT	40.47 53.44 41.01 53.545 ;
		RECT	40.47 53.935 41.01 54.025 ;
		RECT	40.47 54.435 41.01 54.515 ;
		RECT	40.47 54.615 41.01 54.825 ;
		RECT	40.47 54.925 41.01 55.02 ;
		RECT	40.47 55.41 41.01 55.51 ;
		RECT	40.47 55.9 41.01 56.005 ;
		RECT	40.47 56.395 41.01 56.485 ;
		RECT	40.47 56.895 41.01 56.985 ;
		RECT	40.47 57.375 41.01 57.48 ;
		RECT	40.47 57.87 41.01 57.97 ;
		RECT	40.47 58.36 41.01 58.465 ;
		RECT	40.47 58.565 41.01 58.755 ;
		RECT	40.47 58.855 41.01 58.955 ;
		RECT	40.47 59.345 41.01 59.445 ;
		RECT	40.47 59.835 41.01 59.94 ;
		RECT	40.47 60.33 41.01 60.43 ;
		RECT	40.47 60.82 41.01 60.925 ;
		RECT	40.47 61.315 41.01 61.415 ;
		RECT	40.47 61.805 41.01 61.905 ;
		RECT	40.47 62.49 41.01 62.7 ;
		RECT	40.47 62.8 41.01 62.89 ;
		RECT	40.47 63.28 41.01 63.375 ;
		RECT	40.47 63.79 41.01 63.86 ;
		RECT	40.47 64.28 41.01 64.35 ;
		RECT	40.47 64.765 41.01 64.825 ;
		RECT	40.47 65.215 41.01 65.35 ;
		RECT	40.47 65.74 41.01 65.81 ;
		RECT	40.47 66.2 41.01 66.35 ;
		RECT	40.47 66.45 41.01 66.64 ;
		RECT	40.47 66.925 41.01 67.115 ;
		RECT	40.47 67.215 41.01 67.32 ;
		RECT	40.47 68.2 41.01 68.305 ;
		RECT	40.47 68.705 41.01 68.915 ;
		RECT	41.01 29.15 41.55 29.34 ;
		RECT	41.01 29.825 41.55 29.925 ;
		RECT	41.01 30.805 41.55 30.91 ;
		RECT	41.01 31.01 41.55 31.2 ;
		RECT	41.01 31.485 41.55 31.675 ;
		RECT	41.01 31.78 41.55 31.93 ;
		RECT	41.01 32.32 41.55 32.385 ;
		RECT	41.01 32.775 41.55 32.88 ;
		RECT	41.01 33.27 41.55 33.37 ;
		RECT	41.01 34.25 41.55 34.355 ;
		RECT	41.01 34.745 41.55 34.845 ;
		RECT	41.01 35.235 41.55 35.34 ;
		RECT	41.01 35.44 41.55 35.63 ;
		RECT	41.01 35.73 41.55 35.83 ;
		RECT	41.01 36.22 41.55 36.325 ;
		RECT	41.01 36.715 41.55 36.815 ;
		RECT	41.01 37.205 41.55 37.305 ;
		RECT	41.01 37.695 41.55 37.8 ;
		RECT	41.01 38.19 41.55 38.29 ;
		RECT	41.01 38.68 41.55 38.78 ;
		RECT	41.01 39.17 41.55 39.275 ;
		RECT	41.01 39.375 41.55 39.565 ;
		RECT	41.01 39.665 41.55 39.765 ;
		RECT	41.01 40.155 41.55 40.26 ;
		RECT	41.01 40.65 41.55 40.75 ;
		RECT	41.01 41.14 41.55 41.23 ;
		RECT	41.01 41.64 41.55 41.735 ;
		RECT	41.01 42.125 41.55 42.225 ;
		RECT	41.01 42.615 41.55 42.72 ;
		RECT	41.01 43.11 41.55 43.2 ;
		RECT	41.01 43.3 41.55 43.51 ;
		RECT	41.01 43.61 41.55 43.705 ;
		RECT	41.01 44.095 41.55 44.2 ;
		RECT	41.01 44.59 41.55 44.685 ;
		RECT	41.01 45.075 41.55 45.18 ;
		RECT	41.01 45.57 41.55 45.655 ;
		RECT	41.01 46.055 41.55 46.265 ;
		RECT	41.01 46.38 41.55 46.57 ;
		RECT	41.01 47.245 41.55 47.435 ;
		RECT	41.01 48.03 41.55 48.13 ;
		RECT	41.01 48.52 41.55 48.62 ;
		RECT	41.01 49.01 41.55 49.115 ;
		RECT	41.01 49.505 41.55 49.605 ;
		RECT	41.01 49.995 41.55 50.1 ;
		RECT	41.01 50.69 41.55 50.88 ;
		RECT	41.01 51.495 41.55 51.685 ;
		RECT	41.01 51.83 41.55 52.04 ;
		RECT	41.01 52.47 41.55 52.555 ;
		RECT	41.01 52.945 41.55 53.05 ;
		RECT	41.01 53.44 41.55 53.545 ;
		RECT	41.01 53.935 41.55 54.025 ;
		RECT	41.01 54.435 41.55 54.515 ;
		RECT	41.01 54.615 41.55 54.825 ;
		RECT	41.01 54.925 41.55 55.02 ;
		RECT	41.01 55.41 41.55 55.51 ;
		RECT	41.01 55.9 41.55 56.005 ;
		RECT	41.01 56.395 41.55 56.485 ;
		RECT	41.01 56.895 41.55 56.985 ;
		RECT	41.01 57.375 41.55 57.48 ;
		RECT	41.01 57.87 41.55 57.97 ;
		RECT	41.01 58.36 41.55 58.465 ;
		RECT	41.01 58.565 41.55 58.755 ;
		RECT	41.01 58.855 41.55 58.955 ;
		RECT	41.01 59.345 41.55 59.445 ;
		RECT	41.01 59.835 41.55 59.94 ;
		RECT	41.01 60.33 41.55 60.43 ;
		RECT	41.01 60.82 41.55 60.925 ;
		RECT	41.01 61.315 41.55 61.415 ;
		RECT	41.01 61.805 41.55 61.905 ;
		RECT	41.01 62.49 41.55 62.7 ;
		RECT	41.01 62.8 41.55 62.89 ;
		RECT	41.01 63.28 41.55 63.375 ;
		RECT	41.01 63.79 41.55 63.86 ;
		RECT	41.01 64.28 41.55 64.35 ;
		RECT	41.01 64.765 41.55 64.825 ;
		RECT	41.01 65.215 41.55 65.35 ;
		RECT	41.01 65.74 41.55 65.81 ;
		RECT	41.01 66.2 41.55 66.35 ;
		RECT	41.01 66.45 41.55 66.64 ;
		RECT	41.01 66.925 41.55 67.115 ;
		RECT	41.01 67.215 41.55 67.32 ;
		RECT	41.01 68.2 41.55 68.305 ;
		RECT	41.01 68.705 41.55 68.915 ;
		RECT	41.55 29.15 42.09 29.34 ;
		RECT	41.55 29.825 42.09 29.925 ;
		RECT	41.55 30.805 42.09 30.91 ;
		RECT	41.55 31.01 42.09 31.2 ;
		RECT	41.55 31.485 42.09 31.675 ;
		RECT	41.55 31.78 42.09 31.93 ;
		RECT	41.55 32.32 42.09 32.385 ;
		RECT	41.55 32.775 42.09 32.88 ;
		RECT	41.55 33.27 42.09 33.37 ;
		RECT	41.55 34.25 42.09 34.355 ;
		RECT	41.55 34.745 42.09 34.845 ;
		RECT	41.55 35.235 42.09 35.34 ;
		RECT	41.55 35.44 42.09 35.63 ;
		RECT	41.55 35.73 42.09 35.83 ;
		RECT	41.55 36.22 42.09 36.325 ;
		RECT	41.55 36.715 42.09 36.815 ;
		RECT	41.55 37.205 42.09 37.305 ;
		RECT	41.55 37.695 42.09 37.8 ;
		RECT	41.55 38.19 42.09 38.29 ;
		RECT	41.55 38.68 42.09 38.78 ;
		RECT	41.55 39.17 42.09 39.275 ;
		RECT	41.55 39.375 42.09 39.565 ;
		RECT	41.55 39.665 42.09 39.765 ;
		RECT	41.55 40.155 42.09 40.26 ;
		RECT	41.55 40.65 42.09 40.75 ;
		RECT	41.55 41.14 42.09 41.23 ;
		RECT	41.55 41.64 42.09 41.735 ;
		RECT	41.55 42.125 42.09 42.225 ;
		RECT	41.55 42.615 42.09 42.72 ;
		RECT	41.55 43.11 42.09 43.2 ;
		RECT	41.55 43.3 42.09 43.51 ;
		RECT	41.55 43.61 42.09 43.705 ;
		RECT	41.55 44.095 42.09 44.2 ;
		RECT	41.55 44.59 42.09 44.685 ;
		RECT	41.55 45.075 42.09 45.18 ;
		RECT	41.55 45.57 42.09 45.655 ;
		RECT	41.55 46.055 42.09 46.265 ;
		RECT	41.55 46.38 42.09 46.57 ;
		RECT	41.55 47.245 42.09 47.435 ;
		RECT	41.55 48.03 42.09 48.13 ;
		RECT	41.55 48.52 42.09 48.62 ;
		RECT	41.55 49.01 42.09 49.115 ;
		RECT	41.55 49.505 42.09 49.605 ;
		RECT	41.55 49.995 42.09 50.1 ;
		RECT	41.55 50.69 42.09 50.88 ;
		RECT	41.55 51.495 42.09 51.685 ;
		RECT	41.55 51.83 42.09 52.04 ;
		RECT	41.55 52.47 42.09 52.555 ;
		RECT	41.55 52.945 42.09 53.05 ;
		RECT	41.55 53.44 42.09 53.545 ;
		RECT	41.55 53.935 42.09 54.025 ;
		RECT	41.55 54.435 42.09 54.515 ;
		RECT	41.55 54.615 42.09 54.825 ;
		RECT	41.55 54.925 42.09 55.02 ;
		RECT	41.55 55.41 42.09 55.51 ;
		RECT	41.55 55.9 42.09 56.005 ;
		RECT	41.55 56.395 42.09 56.485 ;
		RECT	41.55 56.895 42.09 56.985 ;
		RECT	41.55 57.375 42.09 57.48 ;
		RECT	41.55 57.87 42.09 57.97 ;
		RECT	41.55 58.36 42.09 58.465 ;
		RECT	41.55 58.565 42.09 58.755 ;
		RECT	41.55 58.855 42.09 58.955 ;
		RECT	41.55 59.345 42.09 59.445 ;
		RECT	41.55 59.835 42.09 59.94 ;
		RECT	41.55 60.33 42.09 60.43 ;
		RECT	41.55 60.82 42.09 60.925 ;
		RECT	41.55 61.315 42.09 61.415 ;
		RECT	41.55 61.805 42.09 61.905 ;
		RECT	41.55 62.49 42.09 62.7 ;
		RECT	41.55 62.8 42.09 62.89 ;
		RECT	41.55 63.28 42.09 63.375 ;
		RECT	41.55 63.79 42.09 63.86 ;
		RECT	41.55 64.28 42.09 64.35 ;
		RECT	41.55 64.765 42.09 64.825 ;
		RECT	41.55 65.215 42.09 65.35 ;
		RECT	41.55 65.74 42.09 65.81 ;
		RECT	41.55 66.2 42.09 66.35 ;
		RECT	41.55 66.45 42.09 66.64 ;
		RECT	41.55 66.925 42.09 67.115 ;
		RECT	41.55 67.215 42.09 67.32 ;
		RECT	41.55 68.2 42.09 68.305 ;
		RECT	41.55 68.705 42.09 68.915 ;
		RECT	42.09 29.15 42.63 29.34 ;
		RECT	42.09 29.825 42.63 29.925 ;
		RECT	42.09 30.805 42.63 30.91 ;
		RECT	42.09 31.01 42.63 31.2 ;
		RECT	42.09 31.485 42.63 31.675 ;
		RECT	42.09 31.78 42.63 31.93 ;
		RECT	42.09 32.32 42.63 32.385 ;
		RECT	42.09 32.775 42.63 32.88 ;
		RECT	42.09 33.27 42.63 33.37 ;
		RECT	42.09 34.25 42.63 34.355 ;
		RECT	42.09 34.745 42.63 34.845 ;
		RECT	42.09 35.235 42.63 35.34 ;
		RECT	42.09 35.44 42.63 35.63 ;
		RECT	42.09 35.73 42.63 35.83 ;
		RECT	42.09 36.22 42.63 36.325 ;
		RECT	42.09 36.715 42.63 36.815 ;
		RECT	42.09 37.205 42.63 37.305 ;
		RECT	42.09 37.695 42.63 37.8 ;
		RECT	42.09 38.19 42.63 38.29 ;
		RECT	42.09 38.68 42.63 38.78 ;
		RECT	42.09 39.17 42.63 39.275 ;
		RECT	42.09 39.375 42.63 39.565 ;
		RECT	42.09 39.665 42.63 39.765 ;
		RECT	42.09 40.155 42.63 40.26 ;
		RECT	42.09 40.65 42.63 40.75 ;
		RECT	42.09 41.14 42.63 41.23 ;
		RECT	42.09 41.64 42.63 41.735 ;
		RECT	42.09 42.125 42.63 42.225 ;
		RECT	42.09 42.615 42.63 42.72 ;
		RECT	42.09 43.11 42.63 43.2 ;
		RECT	42.09 43.3 42.63 43.51 ;
		RECT	42.09 43.61 42.63 43.705 ;
		RECT	42.09 44.095 42.63 44.2 ;
		RECT	42.09 44.59 42.63 44.685 ;
		RECT	42.09 45.075 42.63 45.18 ;
		RECT	42.09 45.57 42.63 45.655 ;
		RECT	42.09 46.055 42.63 46.265 ;
		RECT	42.09 46.38 42.63 46.57 ;
		RECT	42.09 47.245 42.63 47.435 ;
		RECT	42.09 48.03 42.63 48.13 ;
		RECT	42.09 48.52 42.63 48.62 ;
		RECT	42.09 49.01 42.63 49.115 ;
		RECT	42.09 49.505 42.63 49.605 ;
		RECT	42.09 49.995 42.63 50.1 ;
		RECT	42.09 50.69 42.63 50.88 ;
		RECT	42.09 51.495 42.63 51.685 ;
		RECT	42.09 51.83 42.63 52.04 ;
		RECT	42.09 52.47 42.63 52.555 ;
		RECT	42.09 52.945 42.63 53.05 ;
		RECT	42.09 53.44 42.63 53.545 ;
		RECT	42.09 53.935 42.63 54.025 ;
		RECT	42.09 54.435 42.63 54.515 ;
		RECT	42.09 54.615 42.63 54.825 ;
		RECT	42.09 54.925 42.63 55.02 ;
		RECT	42.09 55.41 42.63 55.51 ;
		RECT	42.09 55.9 42.63 56.005 ;
		RECT	42.09 56.395 42.63 56.485 ;
		RECT	42.09 56.895 42.63 56.985 ;
		RECT	42.09 57.375 42.63 57.48 ;
		RECT	42.09 57.87 42.63 57.97 ;
		RECT	42.09 58.36 42.63 58.465 ;
		RECT	42.09 58.565 42.63 58.755 ;
		RECT	42.09 58.855 42.63 58.955 ;
		RECT	42.09 59.345 42.63 59.445 ;
		RECT	42.09 59.835 42.63 59.94 ;
		RECT	42.09 60.33 42.63 60.43 ;
		RECT	42.09 60.82 42.63 60.925 ;
		RECT	42.09 61.315 42.63 61.415 ;
		RECT	42.09 61.805 42.63 61.905 ;
		RECT	42.09 62.49 42.63 62.7 ;
		RECT	42.09 62.8 42.63 62.89 ;
		RECT	42.09 63.28 42.63 63.375 ;
		RECT	42.09 63.79 42.63 63.86 ;
		RECT	42.09 64.28 42.63 64.35 ;
		RECT	42.09 64.765 42.63 64.825 ;
		RECT	42.09 65.215 42.63 65.35 ;
		RECT	42.09 65.74 42.63 65.81 ;
		RECT	42.09 66.2 42.63 66.35 ;
		RECT	42.09 66.45 42.63 66.64 ;
		RECT	42.09 66.925 42.63 67.115 ;
		RECT	42.09 67.215 42.63 67.32 ;
		RECT	42.09 68.2 42.63 68.305 ;
		RECT	42.09 68.705 42.63 68.915 ;
		RECT	42.63 29.15 43.17 29.34 ;
		RECT	42.63 29.825 43.17 29.925 ;
		RECT	42.63 30.805 43.17 30.91 ;
		RECT	42.63 31.01 43.17 31.2 ;
		RECT	42.63 31.485 43.17 31.675 ;
		RECT	42.63 31.78 43.17 31.93 ;
		RECT	42.63 32.32 43.17 32.385 ;
		RECT	42.63 32.775 43.17 32.88 ;
		RECT	42.63 33.27 43.17 33.37 ;
		RECT	42.63 34.25 43.17 34.355 ;
		RECT	42.63 34.745 43.17 34.845 ;
		RECT	42.63 35.235 43.17 35.34 ;
		RECT	42.63 35.44 43.17 35.63 ;
		RECT	42.63 35.73 43.17 35.83 ;
		RECT	42.63 36.22 43.17 36.325 ;
		RECT	42.63 36.715 43.17 36.815 ;
		RECT	42.63 37.205 43.17 37.305 ;
		RECT	42.63 37.695 43.17 37.8 ;
		RECT	42.63 38.19 43.17 38.29 ;
		RECT	42.63 38.68 43.17 38.78 ;
		RECT	42.63 39.17 43.17 39.275 ;
		RECT	42.63 39.375 43.17 39.565 ;
		RECT	42.63 39.665 43.17 39.765 ;
		RECT	42.63 40.155 43.17 40.26 ;
		RECT	42.63 40.65 43.17 40.75 ;
		RECT	42.63 41.14 43.17 41.23 ;
		RECT	42.63 41.64 43.17 41.735 ;
		RECT	42.63 42.125 43.17 42.225 ;
		RECT	42.63 42.615 43.17 42.72 ;
		RECT	42.63 43.11 43.17 43.2 ;
		RECT	42.63 43.3 43.17 43.51 ;
		RECT	42.63 43.61 43.17 43.705 ;
		RECT	42.63 44.095 43.17 44.2 ;
		RECT	42.63 44.59 43.17 44.685 ;
		RECT	42.63 45.075 43.17 45.18 ;
		RECT	42.63 45.57 43.17 45.655 ;
		RECT	42.63 46.055 43.17 46.265 ;
		RECT	42.63 46.38 43.17 46.57 ;
		RECT	42.63 47.245 43.17 47.435 ;
		RECT	42.63 48.03 43.17 48.13 ;
		RECT	42.63 48.52 43.17 48.62 ;
		RECT	42.63 49.01 43.17 49.115 ;
		RECT	42.63 49.505 43.17 49.605 ;
		RECT	42.63 49.995 43.17 50.1 ;
		RECT	42.63 50.69 43.17 50.88 ;
		RECT	42.63 51.495 43.17 51.685 ;
		RECT	42.63 51.83 43.17 52.04 ;
		RECT	42.63 52.47 43.17 52.555 ;
		RECT	42.63 52.945 43.17 53.05 ;
		RECT	42.63 53.44 43.17 53.545 ;
		RECT	42.63 53.935 43.17 54.025 ;
		RECT	42.63 54.435 43.17 54.515 ;
		RECT	42.63 54.615 43.17 54.825 ;
		RECT	42.63 54.925 43.17 55.02 ;
		RECT	42.63 55.41 43.17 55.51 ;
		RECT	42.63 55.9 43.17 56.005 ;
		RECT	42.63 56.395 43.17 56.485 ;
		RECT	42.63 56.895 43.17 56.985 ;
		RECT	42.63 57.375 43.17 57.48 ;
		RECT	42.63 57.87 43.17 57.97 ;
		RECT	42.63 58.36 43.17 58.465 ;
		RECT	42.63 58.565 43.17 58.755 ;
		RECT	42.63 58.855 43.17 58.955 ;
		RECT	42.63 59.345 43.17 59.445 ;
		RECT	42.63 59.835 43.17 59.94 ;
		RECT	42.63 60.33 43.17 60.43 ;
		RECT	42.63 60.82 43.17 60.925 ;
		RECT	42.63 61.315 43.17 61.415 ;
		RECT	42.63 61.805 43.17 61.905 ;
		RECT	42.63 62.49 43.17 62.7 ;
		RECT	42.63 62.8 43.17 62.89 ;
		RECT	42.63 63.28 43.17 63.375 ;
		RECT	42.63 63.79 43.17 63.86 ;
		RECT	42.63 64.28 43.17 64.35 ;
		RECT	42.63 64.765 43.17 64.825 ;
		RECT	42.63 65.215 43.17 65.35 ;
		RECT	42.63 65.74 43.17 65.81 ;
		RECT	42.63 66.2 43.17 66.35 ;
		RECT	42.63 66.45 43.17 66.64 ;
		RECT	42.63 66.925 43.17 67.115 ;
		RECT	42.63 67.215 43.17 67.32 ;
		RECT	42.63 68.2 43.17 68.305 ;
		RECT	42.63 68.705 43.17 68.915 ;
		RECT	43.17 29.15 43.71 29.34 ;
		RECT	43.17 29.825 43.71 29.925 ;
		RECT	43.17 30.805 43.71 30.91 ;
		RECT	43.17 31.01 43.71 31.2 ;
		RECT	43.17 31.485 43.71 31.675 ;
		RECT	43.17 31.78 43.71 31.93 ;
		RECT	43.17 32.32 43.71 32.385 ;
		RECT	43.17 32.775 43.71 32.88 ;
		RECT	43.17 33.27 43.71 33.37 ;
		RECT	43.17 34.25 43.71 34.355 ;
		RECT	43.17 34.745 43.71 34.845 ;
		RECT	43.17 35.235 43.71 35.34 ;
		RECT	43.17 35.44 43.71 35.63 ;
		RECT	43.17 35.73 43.71 35.83 ;
		RECT	43.17 36.22 43.71 36.325 ;
		RECT	43.17 36.715 43.71 36.815 ;
		RECT	43.17 37.205 43.71 37.305 ;
		RECT	43.17 37.695 43.71 37.8 ;
		RECT	43.17 38.19 43.71 38.29 ;
		RECT	43.17 38.68 43.71 38.78 ;
		RECT	43.17 39.17 43.71 39.275 ;
		RECT	43.17 39.375 43.71 39.565 ;
		RECT	43.17 39.665 43.71 39.765 ;
		RECT	43.17 40.155 43.71 40.26 ;
		RECT	43.17 40.65 43.71 40.75 ;
		RECT	43.17 41.14 43.71 41.23 ;
		RECT	43.17 41.64 43.71 41.735 ;
		RECT	43.17 42.125 43.71 42.225 ;
		RECT	43.17 42.615 43.71 42.72 ;
		RECT	43.17 43.11 43.71 43.2 ;
		RECT	43.17 43.3 43.71 43.51 ;
		RECT	43.17 43.61 43.71 43.705 ;
		RECT	43.17 44.095 43.71 44.2 ;
		RECT	43.17 44.59 43.71 44.685 ;
		RECT	43.17 45.075 43.71 45.18 ;
		RECT	43.17 45.57 43.71 45.655 ;
		RECT	43.17 46.055 43.71 46.265 ;
		RECT	43.17 46.38 43.71 46.57 ;
		RECT	43.17 47.245 43.71 47.435 ;
		RECT	43.17 48.03 43.71 48.13 ;
		RECT	43.17 48.52 43.71 48.62 ;
		RECT	43.17 49.01 43.71 49.115 ;
		RECT	43.17 49.505 43.71 49.605 ;
		RECT	43.17 49.995 43.71 50.1 ;
		RECT	43.17 50.69 43.71 50.88 ;
		RECT	43.17 51.495 43.71 51.685 ;
		RECT	43.17 51.83 43.71 52.04 ;
		RECT	43.17 52.47 43.71 52.555 ;
		RECT	43.17 52.945 43.71 53.05 ;
		RECT	43.17 53.44 43.71 53.545 ;
		RECT	43.17 53.935 43.71 54.025 ;
		RECT	43.17 54.435 43.71 54.515 ;
		RECT	43.17 54.615 43.71 54.825 ;
		RECT	43.17 54.925 43.71 55.02 ;
		RECT	43.17 55.41 43.71 55.51 ;
		RECT	43.17 55.9 43.71 56.005 ;
		RECT	43.17 56.395 43.71 56.485 ;
		RECT	43.17 56.895 43.71 56.985 ;
		RECT	43.17 57.375 43.71 57.48 ;
		RECT	43.17 57.87 43.71 57.97 ;
		RECT	43.17 58.36 43.71 58.465 ;
		RECT	43.17 58.565 43.71 58.755 ;
		RECT	43.17 58.855 43.71 58.955 ;
		RECT	43.17 59.345 43.71 59.445 ;
		RECT	43.17 59.835 43.71 59.94 ;
		RECT	43.17 60.33 43.71 60.43 ;
		RECT	43.17 60.82 43.71 60.925 ;
		RECT	43.17 61.315 43.71 61.415 ;
		RECT	43.17 61.805 43.71 61.905 ;
		RECT	43.17 62.49 43.71 62.7 ;
		RECT	43.17 62.8 43.71 62.89 ;
		RECT	43.17 63.28 43.71 63.375 ;
		RECT	43.17 63.79 43.71 63.86 ;
		RECT	43.17 64.28 43.71 64.35 ;
		RECT	43.17 64.765 43.71 64.825 ;
		RECT	43.17 65.215 43.71 65.35 ;
		RECT	43.17 65.74 43.71 65.81 ;
		RECT	43.17 66.2 43.71 66.35 ;
		RECT	43.17 66.45 43.71 66.64 ;
		RECT	43.17 66.925 43.71 67.115 ;
		RECT	43.17 67.215 43.71 67.32 ;
		RECT	43.17 68.2 43.71 68.305 ;
		RECT	43.17 68.705 43.71 68.915 ;
		RECT	43.71 29.15 44.25 29.34 ;
		RECT	43.71 29.825 44.25 29.925 ;
		RECT	43.71 30.805 44.25 30.91 ;
		RECT	43.71 31.01 44.25 31.2 ;
		RECT	43.71 31.485 44.25 31.675 ;
		RECT	43.71 31.78 44.25 31.93 ;
		RECT	43.71 32.32 44.25 32.385 ;
		RECT	43.71 32.775 44.25 32.88 ;
		RECT	43.71 33.27 44.25 33.37 ;
		RECT	43.71 34.25 44.25 34.355 ;
		RECT	43.71 34.745 44.25 34.845 ;
		RECT	43.71 35.235 44.25 35.34 ;
		RECT	43.71 35.44 44.25 35.63 ;
		RECT	43.71 35.73 44.25 35.83 ;
		RECT	43.71 36.22 44.25 36.325 ;
		RECT	43.71 36.715 44.25 36.815 ;
		RECT	43.71 37.205 44.25 37.305 ;
		RECT	43.71 37.695 44.25 37.8 ;
		RECT	43.71 38.19 44.25 38.29 ;
		RECT	43.71 38.68 44.25 38.78 ;
		RECT	43.71 39.17 44.25 39.275 ;
		RECT	43.71 39.375 44.25 39.565 ;
		RECT	43.71 39.665 44.25 39.765 ;
		RECT	43.71 40.155 44.25 40.26 ;
		RECT	43.71 40.65 44.25 40.75 ;
		RECT	43.71 41.14 44.25 41.23 ;
		RECT	43.71 41.64 44.25 41.735 ;
		RECT	43.71 42.125 44.25 42.225 ;
		RECT	43.71 42.615 44.25 42.72 ;
		RECT	43.71 43.11 44.25 43.2 ;
		RECT	43.71 43.3 44.25 43.51 ;
		RECT	43.71 43.61 44.25 43.705 ;
		RECT	43.71 44.095 44.25 44.2 ;
		RECT	43.71 44.59 44.25 44.685 ;
		RECT	43.71 45.075 44.25 45.18 ;
		RECT	43.71 45.57 44.25 45.655 ;
		RECT	43.71 46.055 44.25 46.265 ;
		RECT	43.71 46.38 44.25 46.57 ;
		RECT	43.71 47.245 44.25 47.435 ;
		RECT	43.71 48.03 44.25 48.13 ;
		RECT	43.71 48.52 44.25 48.62 ;
		RECT	43.71 49.01 44.25 49.115 ;
		RECT	43.71 49.505 44.25 49.605 ;
		RECT	43.71 49.995 44.25 50.1 ;
		RECT	43.71 50.69 44.25 50.88 ;
		RECT	43.71 51.495 44.25 51.685 ;
		RECT	43.71 51.83 44.25 52.04 ;
		RECT	43.71 52.47 44.25 52.555 ;
		RECT	43.71 52.945 44.25 53.05 ;
		RECT	43.71 53.44 44.25 53.545 ;
		RECT	43.71 53.935 44.25 54.025 ;
		RECT	43.71 54.435 44.25 54.515 ;
		RECT	43.71 54.615 44.25 54.825 ;
		RECT	43.71 54.925 44.25 55.02 ;
		RECT	43.71 55.41 44.25 55.51 ;
		RECT	43.71 55.9 44.25 56.005 ;
		RECT	43.71 56.395 44.25 56.485 ;
		RECT	43.71 56.895 44.25 56.985 ;
		RECT	43.71 57.375 44.25 57.48 ;
		RECT	43.71 57.87 44.25 57.97 ;
		RECT	43.71 58.36 44.25 58.465 ;
		RECT	43.71 58.565 44.25 58.755 ;
		RECT	43.71 58.855 44.25 58.955 ;
		RECT	43.71 59.345 44.25 59.445 ;
		RECT	43.71 59.835 44.25 59.94 ;
		RECT	43.71 60.33 44.25 60.43 ;
		RECT	43.71 60.82 44.25 60.925 ;
		RECT	43.71 61.315 44.25 61.415 ;
		RECT	43.71 61.805 44.25 61.905 ;
		RECT	43.71 62.49 44.25 62.7 ;
		RECT	43.71 62.8 44.25 62.89 ;
		RECT	43.71 63.28 44.25 63.375 ;
		RECT	43.71 63.79 44.25 63.86 ;
		RECT	43.71 64.28 44.25 64.35 ;
		RECT	43.71 64.765 44.25 64.825 ;
		RECT	43.71 65.215 44.25 65.35 ;
		RECT	43.71 65.74 44.25 65.81 ;
		RECT	43.71 66.2 44.25 66.35 ;
		RECT	43.71 66.45 44.25 66.64 ;
		RECT	43.71 66.925 44.25 67.115 ;
		RECT	43.71 67.215 44.25 67.32 ;
		RECT	43.71 68.2 44.25 68.305 ;
		RECT	43.71 68.705 44.25 68.915 ;
		RECT	44.25 29.15 44.79 29.34 ;
		RECT	44.25 29.825 44.79 29.925 ;
		RECT	44.25 30.805 44.79 30.91 ;
		RECT	44.25 31.01 44.79 31.2 ;
		RECT	44.25 31.485 44.79 31.675 ;
		RECT	44.25 31.78 44.79 31.93 ;
		RECT	44.25 32.32 44.79 32.385 ;
		RECT	44.25 32.775 44.79 32.88 ;
		RECT	44.25 33.27 44.79 33.37 ;
		RECT	44.25 34.25 44.79 34.355 ;
		RECT	44.25 34.745 44.79 34.845 ;
		RECT	44.25 35.235 44.79 35.34 ;
		RECT	44.25 35.44 44.79 35.63 ;
		RECT	44.25 35.73 44.79 35.83 ;
		RECT	44.25 36.22 44.79 36.325 ;
		RECT	44.25 36.715 44.79 36.815 ;
		RECT	44.25 37.205 44.79 37.305 ;
		RECT	44.25 37.695 44.79 37.8 ;
		RECT	44.25 38.19 44.79 38.29 ;
		RECT	44.25 38.68 44.79 38.78 ;
		RECT	44.25 39.17 44.79 39.275 ;
		RECT	44.25 39.375 44.79 39.565 ;
		RECT	44.25 39.665 44.79 39.765 ;
		RECT	44.25 40.155 44.79 40.26 ;
		RECT	44.25 40.65 44.79 40.75 ;
		RECT	44.25 41.14 44.79 41.23 ;
		RECT	44.25 41.64 44.79 41.735 ;
		RECT	44.25 42.125 44.79 42.225 ;
		RECT	44.25 42.615 44.79 42.72 ;
		RECT	44.25 43.11 44.79 43.2 ;
		RECT	44.25 43.3 44.79 43.51 ;
		RECT	44.25 43.61 44.79 43.705 ;
		RECT	44.25 44.095 44.79 44.2 ;
		RECT	44.25 44.59 44.79 44.685 ;
		RECT	44.25 45.075 44.79 45.18 ;
		RECT	44.25 45.57 44.79 45.655 ;
		RECT	44.25 46.055 44.79 46.265 ;
		RECT	44.25 46.38 44.79 46.57 ;
		RECT	44.25 47.245 44.79 47.435 ;
		RECT	44.25 48.03 44.79 48.13 ;
		RECT	44.25 48.52 44.79 48.62 ;
		RECT	44.25 49.01 44.79 49.115 ;
		RECT	44.25 49.505 44.79 49.605 ;
		RECT	44.25 49.995 44.79 50.1 ;
		RECT	44.25 50.69 44.79 50.88 ;
		RECT	44.25 51.495 44.79 51.685 ;
		RECT	44.25 51.83 44.79 52.04 ;
		RECT	44.25 52.47 44.79 52.555 ;
		RECT	44.25 52.945 44.79 53.05 ;
		RECT	44.25 53.44 44.79 53.545 ;
		RECT	44.25 53.935 44.79 54.025 ;
		RECT	44.25 54.435 44.79 54.515 ;
		RECT	44.25 54.615 44.79 54.825 ;
		RECT	44.25 54.925 44.79 55.02 ;
		RECT	44.25 55.41 44.79 55.51 ;
		RECT	44.25 55.9 44.79 56.005 ;
		RECT	44.25 56.395 44.79 56.485 ;
		RECT	44.25 56.895 44.79 56.985 ;
		RECT	44.25 57.375 44.79 57.48 ;
		RECT	44.25 57.87 44.79 57.97 ;
		RECT	44.25 58.36 44.79 58.465 ;
		RECT	44.25 58.565 44.79 58.755 ;
		RECT	44.25 58.855 44.79 58.955 ;
		RECT	44.25 59.345 44.79 59.445 ;
		RECT	44.25 59.835 44.79 59.94 ;
		RECT	44.25 60.33 44.79 60.43 ;
		RECT	44.25 60.82 44.79 60.925 ;
		RECT	44.25 61.315 44.79 61.415 ;
		RECT	44.25 61.805 44.79 61.905 ;
		RECT	44.25 62.49 44.79 62.7 ;
		RECT	44.25 62.8 44.79 62.89 ;
		RECT	44.25 63.28 44.79 63.375 ;
		RECT	44.25 63.79 44.79 63.86 ;
		RECT	44.25 64.28 44.79 64.35 ;
		RECT	44.25 64.765 44.79 64.825 ;
		RECT	44.25 65.215 44.79 65.35 ;
		RECT	44.25 65.74 44.79 65.81 ;
		RECT	44.25 66.2 44.79 66.35 ;
		RECT	44.25 66.45 44.79 66.64 ;
		RECT	44.25 66.925 44.79 67.115 ;
		RECT	44.25 67.215 44.79 67.32 ;
		RECT	44.25 68.2 44.79 68.305 ;
		RECT	44.25 68.705 44.79 68.915 ;
		RECT	44.79 29.15 45.33 29.34 ;
		RECT	44.79 29.825 45.33 29.925 ;
		RECT	44.79 30.805 45.33 30.91 ;
		RECT	44.79 31.01 45.33 31.2 ;
		RECT	44.79 31.485 45.33 31.675 ;
		RECT	44.79 31.78 45.33 31.93 ;
		RECT	44.79 32.32 45.33 32.385 ;
		RECT	44.79 32.775 45.33 32.88 ;
		RECT	44.79 33.27 45.33 33.37 ;
		RECT	44.79 34.25 45.33 34.355 ;
		RECT	44.79 34.745 45.33 34.845 ;
		RECT	44.79 35.235 45.33 35.34 ;
		RECT	44.79 35.44 45.33 35.63 ;
		RECT	44.79 35.73 45.33 35.83 ;
		RECT	44.79 36.22 45.33 36.325 ;
		RECT	44.79 36.715 45.33 36.815 ;
		RECT	44.79 37.205 45.33 37.305 ;
		RECT	44.79 37.695 45.33 37.8 ;
		RECT	44.79 38.19 45.33 38.29 ;
		RECT	44.79 38.68 45.33 38.78 ;
		RECT	44.79 39.17 45.33 39.275 ;
		RECT	44.79 39.375 45.33 39.565 ;
		RECT	44.79 39.665 45.33 39.765 ;
		RECT	44.79 40.155 45.33 40.26 ;
		RECT	44.79 40.65 45.33 40.75 ;
		RECT	44.79 41.14 45.33 41.23 ;
		RECT	44.79 41.64 45.33 41.735 ;
		RECT	44.79 42.125 45.33 42.225 ;
		RECT	44.79 42.615 45.33 42.72 ;
		RECT	44.79 43.11 45.33 43.2 ;
		RECT	44.79 43.3 45.33 43.51 ;
		RECT	44.79 43.61 45.33 43.705 ;
		RECT	44.79 44.095 45.33 44.2 ;
		RECT	44.79 44.59 45.33 44.685 ;
		RECT	44.79 45.075 45.33 45.18 ;
		RECT	44.79 45.57 45.33 45.655 ;
		RECT	44.79 46.055 45.33 46.265 ;
		RECT	44.79 46.38 45.33 46.57 ;
		RECT	44.79 47.245 45.33 47.435 ;
		RECT	44.79 48.03 45.33 48.13 ;
		RECT	44.79 48.52 45.33 48.62 ;
		RECT	44.79 49.01 45.33 49.115 ;
		RECT	44.79 49.505 45.33 49.605 ;
		RECT	44.79 49.995 45.33 50.1 ;
		RECT	44.79 50.69 45.33 50.88 ;
		RECT	44.79 51.495 45.33 51.685 ;
		RECT	44.79 51.83 45.33 52.04 ;
		RECT	44.79 52.47 45.33 52.555 ;
		RECT	44.79 52.945 45.33 53.05 ;
		RECT	44.79 53.44 45.33 53.545 ;
		RECT	44.79 53.935 45.33 54.025 ;
		RECT	44.79 54.435 45.33 54.515 ;
		RECT	44.79 54.615 45.33 54.825 ;
		RECT	44.79 54.925 45.33 55.02 ;
		RECT	44.79 55.41 45.33 55.51 ;
		RECT	44.79 55.9 45.33 56.005 ;
		RECT	44.79 56.395 45.33 56.485 ;
		RECT	44.79 56.895 45.33 56.985 ;
		RECT	44.79 57.375 45.33 57.48 ;
		RECT	44.79 57.87 45.33 57.97 ;
		RECT	44.79 58.36 45.33 58.465 ;
		RECT	44.79 58.565 45.33 58.755 ;
		RECT	44.79 58.855 45.33 58.955 ;
		RECT	44.79 59.345 45.33 59.445 ;
		RECT	44.79 59.835 45.33 59.94 ;
		RECT	44.79 60.33 45.33 60.43 ;
		RECT	44.79 60.82 45.33 60.925 ;
		RECT	44.79 61.315 45.33 61.415 ;
		RECT	44.79 61.805 45.33 61.905 ;
		RECT	44.79 62.49 45.33 62.7 ;
		RECT	44.79 62.8 45.33 62.89 ;
		RECT	44.79 63.28 45.33 63.375 ;
		RECT	44.79 63.79 45.33 63.86 ;
		RECT	44.79 64.28 45.33 64.35 ;
		RECT	44.79 64.765 45.33 64.825 ;
		RECT	44.79 65.215 45.33 65.35 ;
		RECT	44.79 65.74 45.33 65.81 ;
		RECT	44.79 66.2 45.33 66.35 ;
		RECT	44.79 66.45 45.33 66.64 ;
		RECT	44.79 66.925 45.33 67.115 ;
		RECT	44.79 67.215 45.33 67.32 ;
		RECT	44.79 68.2 45.33 68.305 ;
		RECT	44.79 68.705 45.33 68.915 ;
		RECT	45.33 29.15 45.87 29.34 ;
		RECT	45.33 29.825 45.87 29.925 ;
		RECT	45.33 30.805 45.87 30.91 ;
		RECT	45.33 31.01 45.87 31.2 ;
		RECT	45.33 31.485 45.87 31.675 ;
		RECT	45.33 31.78 45.87 31.93 ;
		RECT	45.33 32.32 45.87 32.385 ;
		RECT	45.33 32.775 45.87 32.88 ;
		RECT	45.33 33.27 45.87 33.37 ;
		RECT	45.33 34.25 45.87 34.355 ;
		RECT	45.33 34.745 45.87 34.845 ;
		RECT	45.33 35.235 45.87 35.34 ;
		RECT	45.33 35.44 45.87 35.63 ;
		RECT	45.33 35.73 45.87 35.83 ;
		RECT	45.33 36.22 45.87 36.325 ;
		RECT	45.33 36.715 45.87 36.815 ;
		RECT	45.33 37.205 45.87 37.305 ;
		RECT	45.33 37.695 45.87 37.8 ;
		RECT	45.33 38.19 45.87 38.29 ;
		RECT	45.33 38.68 45.87 38.78 ;
		RECT	45.33 39.17 45.87 39.275 ;
		RECT	45.33 39.375 45.87 39.565 ;
		RECT	45.33 39.665 45.87 39.765 ;
		RECT	45.33 40.155 45.87 40.26 ;
		RECT	45.33 40.65 45.87 40.75 ;
		RECT	45.33 41.14 45.87 41.23 ;
		RECT	45.33 41.64 45.87 41.735 ;
		RECT	45.33 42.125 45.87 42.225 ;
		RECT	45.33 42.615 45.87 42.72 ;
		RECT	45.33 43.11 45.87 43.2 ;
		RECT	45.33 43.3 45.87 43.51 ;
		RECT	45.33 43.61 45.87 43.705 ;
		RECT	45.33 44.095 45.87 44.2 ;
		RECT	45.33 44.59 45.87 44.685 ;
		RECT	45.33 45.075 45.87 45.18 ;
		RECT	45.33 45.57 45.87 45.655 ;
		RECT	45.33 46.055 45.87 46.265 ;
		RECT	45.33 46.38 45.87 46.57 ;
		RECT	45.33 47.245 45.87 47.435 ;
		RECT	45.33 48.03 45.87 48.13 ;
		RECT	45.33 48.52 45.87 48.62 ;
		RECT	45.33 49.01 45.87 49.115 ;
		RECT	45.33 49.505 45.87 49.605 ;
		RECT	45.33 49.995 45.87 50.1 ;
		RECT	45.33 50.69 45.87 50.88 ;
		RECT	45.33 51.495 45.87 51.685 ;
		RECT	45.33 51.83 45.87 52.04 ;
		RECT	45.33 52.47 45.87 52.555 ;
		RECT	45.33 52.945 45.87 53.05 ;
		RECT	45.33 53.44 45.87 53.545 ;
		RECT	45.33 53.935 45.87 54.025 ;
		RECT	45.33 54.435 45.87 54.515 ;
		RECT	45.33 54.615 45.87 54.825 ;
		RECT	45.33 54.925 45.87 55.02 ;
		RECT	45.33 55.41 45.87 55.51 ;
		RECT	45.33 55.9 45.87 56.005 ;
		RECT	45.33 56.395 45.87 56.485 ;
		RECT	45.33 56.895 45.87 56.985 ;
		RECT	45.33 57.375 45.87 57.48 ;
		RECT	45.33 57.87 45.87 57.97 ;
		RECT	45.33 58.36 45.87 58.465 ;
		RECT	45.33 58.565 45.87 58.755 ;
		RECT	45.33 58.855 45.87 58.955 ;
		RECT	45.33 59.345 45.87 59.445 ;
		RECT	45.33 59.835 45.87 59.94 ;
		RECT	45.33 60.33 45.87 60.43 ;
		RECT	45.33 60.82 45.87 60.925 ;
		RECT	45.33 61.315 45.87 61.415 ;
		RECT	45.33 61.805 45.87 61.905 ;
		RECT	45.33 62.49 45.87 62.7 ;
		RECT	45.33 62.8 45.87 62.89 ;
		RECT	45.33 63.28 45.87 63.375 ;
		RECT	45.33 63.79 45.87 63.86 ;
		RECT	45.33 64.28 45.87 64.35 ;
		RECT	45.33 64.765 45.87 64.825 ;
		RECT	45.33 65.215 45.87 65.35 ;
		RECT	45.33 65.74 45.87 65.81 ;
		RECT	45.33 66.2 45.87 66.35 ;
		RECT	45.33 66.45 45.87 66.64 ;
		RECT	45.33 66.925 45.87 67.115 ;
		RECT	45.33 67.215 45.87 67.32 ;
		RECT	45.33 68.2 45.87 68.305 ;
		RECT	45.33 68.705 45.87 68.915 ;
		RECT	45.87 29.15 46.41 29.34 ;
		RECT	45.87 29.825 46.41 29.925 ;
		RECT	45.87 30.805 46.41 30.91 ;
		RECT	45.87 31.01 46.41 31.2 ;
		RECT	45.87 31.485 46.41 31.675 ;
		RECT	45.87 31.78 46.41 31.93 ;
		RECT	45.87 32.32 46.41 32.385 ;
		RECT	45.87 32.775 46.41 32.88 ;
		RECT	45.87 33.27 46.41 33.37 ;
		RECT	45.87 34.25 46.41 34.355 ;
		RECT	45.87 34.745 46.41 34.845 ;
		RECT	45.87 35.235 46.41 35.34 ;
		RECT	45.87 35.44 46.41 35.63 ;
		RECT	45.87 35.73 46.41 35.83 ;
		RECT	45.87 36.22 46.41 36.325 ;
		RECT	45.87 36.715 46.41 36.815 ;
		RECT	45.87 37.205 46.41 37.305 ;
		RECT	45.87 37.695 46.41 37.8 ;
		RECT	45.87 38.19 46.41 38.29 ;
		RECT	45.87 38.68 46.41 38.78 ;
		RECT	45.87 39.17 46.41 39.275 ;
		RECT	45.87 39.375 46.41 39.565 ;
		RECT	45.87 39.665 46.41 39.765 ;
		RECT	45.87 40.155 46.41 40.26 ;
		RECT	45.87 40.65 46.41 40.75 ;
		RECT	45.87 41.14 46.41 41.23 ;
		RECT	45.87 41.64 46.41 41.735 ;
		RECT	45.87 42.125 46.41 42.225 ;
		RECT	45.87 42.615 46.41 42.72 ;
		RECT	45.87 43.11 46.41 43.2 ;
		RECT	45.87 43.3 46.41 43.51 ;
		RECT	45.87 43.61 46.41 43.705 ;
		RECT	45.87 44.095 46.41 44.2 ;
		RECT	45.87 44.59 46.41 44.685 ;
		RECT	45.87 45.075 46.41 45.18 ;
		RECT	45.87 45.57 46.41 45.655 ;
		RECT	45.87 46.055 46.41 46.265 ;
		RECT	45.87 46.38 46.41 46.57 ;
		RECT	45.87 47.245 46.41 47.435 ;
		RECT	45.87 48.03 46.41 48.13 ;
		RECT	45.87 48.52 46.41 48.62 ;
		RECT	45.87 49.01 46.41 49.115 ;
		RECT	45.87 49.505 46.41 49.605 ;
		RECT	45.87 49.995 46.41 50.1 ;
		RECT	45.87 50.69 46.41 50.88 ;
		RECT	45.87 51.495 46.41 51.685 ;
		RECT	45.87 51.83 46.41 52.04 ;
		RECT	45.87 52.47 46.41 52.555 ;
		RECT	45.87 52.945 46.41 53.05 ;
		RECT	45.87 53.44 46.41 53.545 ;
		RECT	45.87 53.935 46.41 54.025 ;
		RECT	45.87 54.435 46.41 54.515 ;
		RECT	45.87 54.615 46.41 54.825 ;
		RECT	45.87 54.925 46.41 55.02 ;
		RECT	45.87 55.41 46.41 55.51 ;
		RECT	45.87 55.9 46.41 56.005 ;
		RECT	45.87 56.395 46.41 56.485 ;
		RECT	45.87 56.895 46.41 56.985 ;
		RECT	45.87 57.375 46.41 57.48 ;
		RECT	45.87 57.87 46.41 57.97 ;
		RECT	45.87 58.36 46.41 58.465 ;
		RECT	45.87 58.565 46.41 58.755 ;
		RECT	45.87 58.855 46.41 58.955 ;
		RECT	45.87 59.345 46.41 59.445 ;
		RECT	45.87 59.835 46.41 59.94 ;
		RECT	45.87 60.33 46.41 60.43 ;
		RECT	45.87 60.82 46.41 60.925 ;
		RECT	45.87 61.315 46.41 61.415 ;
		RECT	45.87 61.805 46.41 61.905 ;
		RECT	45.87 62.49 46.41 62.7 ;
		RECT	45.87 62.8 46.41 62.89 ;
		RECT	45.87 63.28 46.41 63.375 ;
		RECT	45.87 63.79 46.41 63.86 ;
		RECT	45.87 64.28 46.41 64.35 ;
		RECT	45.87 64.765 46.41 64.825 ;
		RECT	45.87 65.215 46.41 65.35 ;
		RECT	45.87 65.74 46.41 65.81 ;
		RECT	45.87 66.2 46.41 66.35 ;
		RECT	45.87 66.45 46.41 66.64 ;
		RECT	45.87 66.925 46.41 67.115 ;
		RECT	45.87 67.215 46.41 67.32 ;
		RECT	45.87 68.2 46.41 68.305 ;
		RECT	45.87 68.705 46.41 68.915 ;
		RECT	46.41 29.15 46.95 29.34 ;
		RECT	46.41 29.825 46.95 29.925 ;
		RECT	46.41 30.805 46.95 30.91 ;
		RECT	46.41 31.01 46.95 31.2 ;
		RECT	46.41 31.485 46.95 31.675 ;
		RECT	46.41 31.78 46.95 31.93 ;
		RECT	46.41 32.32 46.95 32.385 ;
		RECT	46.41 32.775 46.95 32.88 ;
		RECT	46.41 33.27 46.95 33.37 ;
		RECT	46.41 34.25 46.95 34.355 ;
		RECT	46.41 34.745 46.95 34.845 ;
		RECT	46.41 35.235 46.95 35.34 ;
		RECT	46.41 35.44 46.95 35.63 ;
		RECT	46.41 35.73 46.95 35.83 ;
		RECT	46.41 36.22 46.95 36.325 ;
		RECT	46.41 36.715 46.95 36.815 ;
		RECT	46.41 37.205 46.95 37.305 ;
		RECT	46.41 37.695 46.95 37.8 ;
		RECT	46.41 38.19 46.95 38.29 ;
		RECT	46.41 38.68 46.95 38.78 ;
		RECT	46.41 39.17 46.95 39.275 ;
		RECT	46.41 39.375 46.95 39.565 ;
		RECT	46.41 39.665 46.95 39.765 ;
		RECT	46.41 40.155 46.95 40.26 ;
		RECT	46.41 40.65 46.95 40.75 ;
		RECT	46.41 41.14 46.95 41.23 ;
		RECT	46.41 41.64 46.95 41.735 ;
		RECT	46.41 42.125 46.95 42.225 ;
		RECT	46.41 42.615 46.95 42.72 ;
		RECT	46.41 43.11 46.95 43.2 ;
		RECT	46.41 43.3 46.95 43.51 ;
		RECT	46.41 43.61 46.95 43.705 ;
		RECT	46.41 44.095 46.95 44.2 ;
		RECT	46.41 44.59 46.95 44.685 ;
		RECT	46.41 45.075 46.95 45.18 ;
		RECT	46.41 45.57 46.95 45.655 ;
		RECT	46.41 46.055 46.95 46.265 ;
		RECT	46.41 46.38 46.95 46.57 ;
		RECT	46.41 47.245 46.95 47.435 ;
		RECT	46.41 48.03 46.95 48.13 ;
		RECT	46.41 48.52 46.95 48.62 ;
		RECT	46.41 49.01 46.95 49.115 ;
		RECT	46.41 49.505 46.95 49.605 ;
		RECT	46.41 49.995 46.95 50.1 ;
		RECT	46.41 50.69 46.95 50.88 ;
		RECT	46.41 51.495 46.95 51.685 ;
		RECT	46.41 51.83 46.95 52.04 ;
		RECT	46.41 52.47 46.95 52.555 ;
		RECT	46.41 52.945 46.95 53.05 ;
		RECT	46.41 53.44 46.95 53.545 ;
		RECT	46.41 53.935 46.95 54.025 ;
		RECT	46.41 54.435 46.95 54.515 ;
		RECT	46.41 54.615 46.95 54.825 ;
		RECT	46.41 54.925 46.95 55.02 ;
		RECT	46.41 55.41 46.95 55.51 ;
		RECT	46.41 55.9 46.95 56.005 ;
		RECT	46.41 56.395 46.95 56.485 ;
		RECT	46.41 56.895 46.95 56.985 ;
		RECT	46.41 57.375 46.95 57.48 ;
		RECT	46.41 57.87 46.95 57.97 ;
		RECT	46.41 58.36 46.95 58.465 ;
		RECT	46.41 58.565 46.95 58.755 ;
		RECT	46.41 58.855 46.95 58.955 ;
		RECT	46.41 59.345 46.95 59.445 ;
		RECT	46.41 59.835 46.95 59.94 ;
		RECT	46.41 60.33 46.95 60.43 ;
		RECT	46.41 60.82 46.95 60.925 ;
		RECT	46.41 61.315 46.95 61.415 ;
		RECT	46.41 61.805 46.95 61.905 ;
		RECT	46.41 62.49 46.95 62.7 ;
		RECT	46.41 62.8 46.95 62.89 ;
		RECT	46.41 63.28 46.95 63.375 ;
		RECT	46.41 63.79 46.95 63.86 ;
		RECT	46.41 64.28 46.95 64.35 ;
		RECT	46.41 64.765 46.95 64.825 ;
		RECT	46.41 65.215 46.95 65.35 ;
		RECT	46.41 65.74 46.95 65.81 ;
		RECT	46.41 66.2 46.95 66.35 ;
		RECT	46.41 66.45 46.95 66.64 ;
		RECT	46.41 66.925 46.95 67.115 ;
		RECT	46.41 67.215 46.95 67.32 ;
		RECT	46.41 68.2 46.95 68.305 ;
		RECT	46.41 68.705 46.95 68.915 ;
		RECT	46.95 29.15 47.49 29.34 ;
		RECT	46.95 29.825 47.49 29.925 ;
		RECT	46.95 30.805 47.49 30.91 ;
		RECT	46.95 31.01 47.49 31.2 ;
		RECT	46.95 31.485 47.49 31.675 ;
		RECT	46.95 31.78 47.49 31.93 ;
		RECT	46.95 32.32 47.49 32.385 ;
		RECT	46.95 32.775 47.49 32.88 ;
		RECT	46.95 33.27 47.49 33.37 ;
		RECT	46.95 34.25 47.49 34.355 ;
		RECT	46.95 34.745 47.49 34.845 ;
		RECT	46.95 35.235 47.49 35.34 ;
		RECT	46.95 35.44 47.49 35.63 ;
		RECT	46.95 35.73 47.49 35.83 ;
		RECT	46.95 36.22 47.49 36.325 ;
		RECT	46.95 36.715 47.49 36.815 ;
		RECT	46.95 37.205 47.49 37.305 ;
		RECT	46.95 37.695 47.49 37.8 ;
		RECT	46.95 38.19 47.49 38.29 ;
		RECT	46.95 38.68 47.49 38.78 ;
		RECT	46.95 39.17 47.49 39.275 ;
		RECT	46.95 39.375 47.49 39.565 ;
		RECT	46.95 39.665 47.49 39.765 ;
		RECT	46.95 40.155 47.49 40.26 ;
		RECT	46.95 40.65 47.49 40.75 ;
		RECT	46.95 41.14 47.49 41.23 ;
		RECT	46.95 41.64 47.49 41.735 ;
		RECT	46.95 42.125 47.49 42.225 ;
		RECT	46.95 42.615 47.49 42.72 ;
		RECT	46.95 43.11 47.49 43.2 ;
		RECT	46.95 43.3 47.49 43.51 ;
		RECT	46.95 43.61 47.49 43.705 ;
		RECT	46.95 44.095 47.49 44.2 ;
		RECT	46.95 44.59 47.49 44.685 ;
		RECT	46.95 45.075 47.49 45.18 ;
		RECT	46.95 45.57 47.49 45.655 ;
		RECT	46.95 46.055 47.49 46.265 ;
		RECT	46.95 46.38 47.49 46.57 ;
		RECT	46.95 47.245 47.49 47.435 ;
		RECT	46.95 48.03 47.49 48.13 ;
		RECT	46.95 48.52 47.49 48.62 ;
		RECT	46.95 49.01 47.49 49.115 ;
		RECT	46.95 49.505 47.49 49.605 ;
		RECT	46.95 49.995 47.49 50.1 ;
		RECT	46.95 50.69 47.49 50.88 ;
		RECT	46.95 51.495 47.49 51.685 ;
		RECT	46.95 51.83 47.49 52.04 ;
		RECT	46.95 52.47 47.49 52.555 ;
		RECT	46.95 52.945 47.49 53.05 ;
		RECT	46.95 53.44 47.49 53.545 ;
		RECT	46.95 53.935 47.49 54.025 ;
		RECT	46.95 54.435 47.49 54.515 ;
		RECT	46.95 54.615 47.49 54.825 ;
		RECT	46.95 54.925 47.49 55.02 ;
		RECT	46.95 55.41 47.49 55.51 ;
		RECT	46.95 55.9 47.49 56.005 ;
		RECT	46.95 56.395 47.49 56.485 ;
		RECT	46.95 56.895 47.49 56.985 ;
		RECT	46.95 57.375 47.49 57.48 ;
		RECT	46.95 57.87 47.49 57.97 ;
		RECT	46.95 58.36 47.49 58.465 ;
		RECT	46.95 58.565 47.49 58.755 ;
		RECT	46.95 58.855 47.49 58.955 ;
		RECT	46.95 59.345 47.49 59.445 ;
		RECT	46.95 59.835 47.49 59.94 ;
		RECT	46.95 60.33 47.49 60.43 ;
		RECT	46.95 60.82 47.49 60.925 ;
		RECT	46.95 61.315 47.49 61.415 ;
		RECT	46.95 61.805 47.49 61.905 ;
		RECT	46.95 62.49 47.49 62.7 ;
		RECT	46.95 62.8 47.49 62.89 ;
		RECT	46.95 63.28 47.49 63.375 ;
		RECT	46.95 63.79 47.49 63.86 ;
		RECT	46.95 64.28 47.49 64.35 ;
		RECT	46.95 64.765 47.49 64.825 ;
		RECT	46.95 65.215 47.49 65.35 ;
		RECT	46.95 65.74 47.49 65.81 ;
		RECT	46.95 66.2 47.49 66.35 ;
		RECT	46.95 66.45 47.49 66.64 ;
		RECT	46.95 66.925 47.49 67.115 ;
		RECT	46.95 67.215 47.49 67.32 ;
		RECT	46.95 68.2 47.49 68.305 ;
		RECT	46.95 68.705 47.49 68.915 ;
		RECT	47.49 29.15 48.03 29.34 ;
		RECT	47.49 29.825 48.03 29.925 ;
		RECT	47.49 30.805 48.03 30.91 ;
		RECT	47.49 31.01 48.03 31.2 ;
		RECT	47.49 31.485 48.03 31.675 ;
		RECT	47.49 31.78 48.03 31.93 ;
		RECT	47.49 32.32 48.03 32.385 ;
		RECT	47.49 32.775 48.03 32.88 ;
		RECT	47.49 33.27 48.03 33.37 ;
		RECT	47.49 34.25 48.03 34.355 ;
		RECT	47.49 34.745 48.03 34.845 ;
		RECT	47.49 35.235 48.03 35.34 ;
		RECT	47.49 35.44 48.03 35.63 ;
		RECT	47.49 35.73 48.03 35.83 ;
		RECT	47.49 36.22 48.03 36.325 ;
		RECT	47.49 36.715 48.03 36.815 ;
		RECT	47.49 37.205 48.03 37.305 ;
		RECT	47.49 37.695 48.03 37.8 ;
		RECT	47.49 38.19 48.03 38.29 ;
		RECT	47.49 38.68 48.03 38.78 ;
		RECT	47.49 39.17 48.03 39.275 ;
		RECT	47.49 39.375 48.03 39.565 ;
		RECT	47.49 39.665 48.03 39.765 ;
		RECT	47.49 40.155 48.03 40.26 ;
		RECT	47.49 40.65 48.03 40.75 ;
		RECT	47.49 41.14 48.03 41.23 ;
		RECT	47.49 41.64 48.03 41.735 ;
		RECT	47.49 42.125 48.03 42.225 ;
		RECT	47.49 42.615 48.03 42.72 ;
		RECT	47.49 43.11 48.03 43.2 ;
		RECT	47.49 43.3 48.03 43.51 ;
		RECT	47.49 43.61 48.03 43.705 ;
		RECT	47.49 44.095 48.03 44.2 ;
		RECT	47.49 44.59 48.03 44.685 ;
		RECT	47.49 45.075 48.03 45.18 ;
		RECT	47.49 45.57 48.03 45.655 ;
		RECT	47.49 46.055 48.03 46.265 ;
		RECT	47.49 46.38 48.03 46.57 ;
		RECT	47.49 47.245 48.03 47.435 ;
		RECT	47.49 48.03 48.03 48.13 ;
		RECT	47.49 48.52 48.03 48.62 ;
		RECT	47.49 49.01 48.03 49.115 ;
		RECT	47.49 49.505 48.03 49.605 ;
		RECT	47.49 49.995 48.03 50.1 ;
		RECT	47.49 50.69 48.03 50.88 ;
		RECT	47.49 51.495 48.03 51.685 ;
		RECT	47.49 51.83 48.03 52.04 ;
		RECT	47.49 52.47 48.03 52.555 ;
		RECT	47.49 52.945 48.03 53.05 ;
		RECT	47.49 53.44 48.03 53.545 ;
		RECT	47.49 53.935 48.03 54.025 ;
		RECT	47.49 54.435 48.03 54.515 ;
		RECT	47.49 54.615 48.03 54.825 ;
		RECT	47.49 54.925 48.03 55.02 ;
		RECT	47.49 55.41 48.03 55.51 ;
		RECT	47.49 55.9 48.03 56.005 ;
		RECT	47.49 56.395 48.03 56.485 ;
		RECT	47.49 56.895 48.03 56.985 ;
		RECT	47.49 57.375 48.03 57.48 ;
		RECT	47.49 57.87 48.03 57.97 ;
		RECT	47.49 58.36 48.03 58.465 ;
		RECT	47.49 58.565 48.03 58.755 ;
		RECT	47.49 58.855 48.03 58.955 ;
		RECT	47.49 59.345 48.03 59.445 ;
		RECT	47.49 59.835 48.03 59.94 ;
		RECT	47.49 60.33 48.03 60.43 ;
		RECT	47.49 60.82 48.03 60.925 ;
		RECT	47.49 61.315 48.03 61.415 ;
		RECT	47.49 61.805 48.03 61.905 ;
		RECT	47.49 62.49 48.03 62.7 ;
		RECT	47.49 62.8 48.03 62.89 ;
		RECT	47.49 63.28 48.03 63.375 ;
		RECT	47.49 63.79 48.03 63.86 ;
		RECT	47.49 64.28 48.03 64.35 ;
		RECT	47.49 64.765 48.03 64.825 ;
		RECT	47.49 65.215 48.03 65.35 ;
		RECT	47.49 65.74 48.03 65.81 ;
		RECT	47.49 66.2 48.03 66.35 ;
		RECT	47.49 66.45 48.03 66.64 ;
		RECT	47.49 66.925 48.03 67.115 ;
		RECT	47.49 67.215 48.03 67.32 ;
		RECT	47.49 68.2 48.03 68.305 ;
		RECT	47.49 68.705 48.03 68.915 ;
		RECT	48.03 29.15 48.57 29.34 ;
		RECT	48.03 29.825 48.57 29.925 ;
		RECT	48.03 30.805 48.57 30.91 ;
		RECT	48.03 31.01 48.57 31.2 ;
		RECT	48.03 31.485 48.57 31.675 ;
		RECT	48.03 31.78 48.57 31.93 ;
		RECT	48.03 32.32 48.57 32.385 ;
		RECT	48.03 32.775 48.57 32.88 ;
		RECT	48.03 33.27 48.57 33.37 ;
		RECT	48.03 34.25 48.57 34.355 ;
		RECT	48.03 34.745 48.57 34.845 ;
		RECT	48.03 35.235 48.57 35.34 ;
		RECT	48.03 35.44 48.57 35.63 ;
		RECT	48.03 35.73 48.57 35.83 ;
		RECT	48.03 36.22 48.57 36.325 ;
		RECT	48.03 36.715 48.57 36.815 ;
		RECT	48.03 37.205 48.57 37.305 ;
		RECT	48.03 37.695 48.57 37.8 ;
		RECT	48.03 38.19 48.57 38.29 ;
		RECT	48.03 38.68 48.57 38.78 ;
		RECT	48.03 39.17 48.57 39.275 ;
		RECT	48.03 39.375 48.57 39.565 ;
		RECT	48.03 39.665 48.57 39.765 ;
		RECT	48.03 40.155 48.57 40.26 ;
		RECT	48.03 40.65 48.57 40.75 ;
		RECT	48.03 41.14 48.57 41.23 ;
		RECT	48.03 41.64 48.57 41.735 ;
		RECT	48.03 42.125 48.57 42.225 ;
		RECT	48.03 42.615 48.57 42.72 ;
		RECT	48.03 43.11 48.57 43.2 ;
		RECT	48.03 43.3 48.57 43.51 ;
		RECT	48.03 43.61 48.57 43.705 ;
		RECT	48.03 44.095 48.57 44.2 ;
		RECT	48.03 44.59 48.57 44.685 ;
		RECT	48.03 45.075 48.57 45.18 ;
		RECT	48.03 45.57 48.57 45.655 ;
		RECT	48.03 46.055 48.57 46.265 ;
		RECT	48.03 46.38 48.57 46.57 ;
		RECT	48.03 47.245 48.57 47.435 ;
		RECT	48.03 48.03 48.57 48.13 ;
		RECT	48.03 48.52 48.57 48.62 ;
		RECT	48.03 49.01 48.57 49.115 ;
		RECT	48.03 49.505 48.57 49.605 ;
		RECT	48.03 49.995 48.57 50.1 ;
		RECT	48.03 50.69 48.57 50.88 ;
		RECT	48.03 51.495 48.57 51.685 ;
		RECT	48.03 51.83 48.57 52.04 ;
		RECT	48.03 52.47 48.57 52.555 ;
		RECT	48.03 52.945 48.57 53.05 ;
		RECT	48.03 53.44 48.57 53.545 ;
		RECT	48.03 53.935 48.57 54.025 ;
		RECT	48.03 54.435 48.57 54.515 ;
		RECT	48.03 54.615 48.57 54.825 ;
		RECT	48.03 54.925 48.57 55.02 ;
		RECT	48.03 55.41 48.57 55.51 ;
		RECT	48.03 55.9 48.57 56.005 ;
		RECT	48.03 56.395 48.57 56.485 ;
		RECT	48.03 56.895 48.57 56.985 ;
		RECT	48.03 57.375 48.57 57.48 ;
		RECT	48.03 57.87 48.57 57.97 ;
		RECT	48.03 58.36 48.57 58.465 ;
		RECT	48.03 58.565 48.57 58.755 ;
		RECT	48.03 58.855 48.57 58.955 ;
		RECT	48.03 59.345 48.57 59.445 ;
		RECT	48.03 59.835 48.57 59.94 ;
		RECT	48.03 60.33 48.57 60.43 ;
		RECT	48.03 60.82 48.57 60.925 ;
		RECT	48.03 61.315 48.57 61.415 ;
		RECT	48.03 61.805 48.57 61.905 ;
		RECT	48.03 62.49 48.57 62.7 ;
		RECT	48.03 62.8 48.57 62.89 ;
		RECT	48.03 63.28 48.57 63.375 ;
		RECT	48.03 63.79 48.57 63.86 ;
		RECT	48.03 64.28 48.57 64.35 ;
		RECT	48.03 64.765 48.57 64.825 ;
		RECT	48.03 65.215 48.57 65.35 ;
		RECT	48.03 65.74 48.57 65.81 ;
		RECT	48.03 66.2 48.57 66.35 ;
		RECT	48.03 66.45 48.57 66.64 ;
		RECT	48.03 66.925 48.57 67.115 ;
		RECT	48.03 67.215 48.57 67.32 ;
		RECT	48.03 68.2 48.57 68.305 ;
		RECT	48.03 68.705 48.57 68.915 ;
		RECT	48.57 29.15 49.11 29.34 ;
		RECT	48.57 29.825 49.11 29.925 ;
		RECT	48.57 30.805 49.11 30.91 ;
		RECT	48.57 31.01 49.11 31.2 ;
		RECT	48.57 31.485 49.11 31.675 ;
		RECT	48.57 31.78 49.11 31.93 ;
		RECT	48.57 32.32 49.11 32.385 ;
		RECT	48.57 32.775 49.11 32.88 ;
		RECT	48.57 33.27 49.11 33.37 ;
		RECT	48.57 34.25 49.11 34.355 ;
		RECT	48.57 34.745 49.11 34.845 ;
		RECT	48.57 35.235 49.11 35.34 ;
		RECT	48.57 35.44 49.11 35.63 ;
		RECT	48.57 35.73 49.11 35.83 ;
		RECT	48.57 36.22 49.11 36.325 ;
		RECT	48.57 36.715 49.11 36.815 ;
		RECT	48.57 37.205 49.11 37.305 ;
		RECT	48.57 37.695 49.11 37.8 ;
		RECT	48.57 38.19 49.11 38.29 ;
		RECT	48.57 38.68 49.11 38.78 ;
		RECT	48.57 39.17 49.11 39.275 ;
		RECT	48.57 39.375 49.11 39.565 ;
		RECT	48.57 39.665 49.11 39.765 ;
		RECT	48.57 40.155 49.11 40.26 ;
		RECT	48.57 40.65 49.11 40.75 ;
		RECT	48.57 41.14 49.11 41.23 ;
		RECT	48.57 41.64 49.11 41.735 ;
		RECT	48.57 42.125 49.11 42.225 ;
		RECT	48.57 42.615 49.11 42.72 ;
		RECT	48.57 43.11 49.11 43.2 ;
		RECT	48.57 43.3 49.11 43.51 ;
		RECT	48.57 43.61 49.11 43.705 ;
		RECT	48.57 44.095 49.11 44.2 ;
		RECT	48.57 44.59 49.11 44.685 ;
		RECT	48.57 45.075 49.11 45.18 ;
		RECT	48.57 45.57 49.11 45.655 ;
		RECT	48.57 46.055 49.11 46.265 ;
		RECT	48.57 46.38 49.11 46.57 ;
		RECT	48.57 47.245 49.11 47.435 ;
		RECT	48.57 48.03 49.11 48.13 ;
		RECT	48.57 48.52 49.11 48.62 ;
		RECT	48.57 49.01 49.11 49.115 ;
		RECT	48.57 49.505 49.11 49.605 ;
		RECT	48.57 49.995 49.11 50.1 ;
		RECT	48.57 50.69 49.11 50.88 ;
		RECT	48.57 51.495 49.11 51.685 ;
		RECT	48.57 51.83 49.11 52.04 ;
		RECT	48.57 52.47 49.11 52.555 ;
		RECT	48.57 52.945 49.11 53.05 ;
		RECT	48.57 53.44 49.11 53.545 ;
		RECT	48.57 53.935 49.11 54.025 ;
		RECT	48.57 54.435 49.11 54.515 ;
		RECT	48.57 54.615 49.11 54.825 ;
		RECT	48.57 54.925 49.11 55.02 ;
		RECT	48.57 55.41 49.11 55.51 ;
		RECT	48.57 55.9 49.11 56.005 ;
		RECT	48.57 56.395 49.11 56.485 ;
		RECT	48.57 56.895 49.11 56.985 ;
		RECT	48.57 57.375 49.11 57.48 ;
		RECT	48.57 57.87 49.11 57.97 ;
		RECT	48.57 58.36 49.11 58.465 ;
		RECT	48.57 58.565 49.11 58.755 ;
		RECT	48.57 58.855 49.11 58.955 ;
		RECT	48.57 59.345 49.11 59.445 ;
		RECT	48.57 59.835 49.11 59.94 ;
		RECT	48.57 60.33 49.11 60.43 ;
		RECT	48.57 60.82 49.11 60.925 ;
		RECT	48.57 61.315 49.11 61.415 ;
		RECT	48.57 61.805 49.11 61.905 ;
		RECT	48.57 62.49 49.11 62.7 ;
		RECT	48.57 62.8 49.11 62.89 ;
		RECT	48.57 63.28 49.11 63.375 ;
		RECT	48.57 63.79 49.11 63.86 ;
		RECT	48.57 64.28 49.11 64.35 ;
		RECT	48.57 64.765 49.11 64.825 ;
		RECT	48.57 65.215 49.11 65.35 ;
		RECT	48.57 65.74 49.11 65.81 ;
		RECT	48.57 66.2 49.11 66.35 ;
		RECT	48.57 66.45 49.11 66.64 ;
		RECT	48.57 66.925 49.11 67.115 ;
		RECT	48.57 67.215 49.11 67.32 ;
		RECT	48.57 68.2 49.11 68.305 ;
		RECT	48.57 68.705 49.11 68.915 ;
		RECT	49.11 29.15 49.65 29.34 ;
		RECT	49.11 29.825 49.65 29.925 ;
		RECT	49.11 30.805 49.65 30.91 ;
		RECT	49.11 31.01 49.65 31.2 ;
		RECT	49.11 31.485 49.65 31.675 ;
		RECT	49.11 31.78 49.65 31.93 ;
		RECT	49.11 32.32 49.65 32.385 ;
		RECT	49.11 32.775 49.65 32.88 ;
		RECT	49.11 33.27 49.65 33.37 ;
		RECT	49.11 34.25 49.65 34.355 ;
		RECT	49.11 34.745 49.65 34.845 ;
		RECT	49.11 35.235 49.65 35.34 ;
		RECT	49.11 35.44 49.65 35.63 ;
		RECT	49.11 35.73 49.65 35.83 ;
		RECT	49.11 36.22 49.65 36.325 ;
		RECT	49.11 36.715 49.65 36.815 ;
		RECT	49.11 37.205 49.65 37.305 ;
		RECT	49.11 37.695 49.65 37.8 ;
		RECT	49.11 38.19 49.65 38.29 ;
		RECT	49.11 38.68 49.65 38.78 ;
		RECT	49.11 39.17 49.65 39.275 ;
		RECT	49.11 39.375 49.65 39.565 ;
		RECT	49.11 39.665 49.65 39.765 ;
		RECT	49.11 40.155 49.65 40.26 ;
		RECT	49.11 40.65 49.65 40.75 ;
		RECT	49.11 41.14 49.65 41.23 ;
		RECT	49.11 41.64 49.65 41.735 ;
		RECT	49.11 42.125 49.65 42.225 ;
		RECT	49.11 42.615 49.65 42.72 ;
		RECT	49.11 43.11 49.65 43.2 ;
		RECT	49.11 43.3 49.65 43.51 ;
		RECT	49.11 43.61 49.65 43.705 ;
		RECT	49.11 44.095 49.65 44.2 ;
		RECT	49.11 44.59 49.65 44.685 ;
		RECT	49.11 45.075 49.65 45.18 ;
		RECT	49.11 45.57 49.65 45.655 ;
		RECT	49.11 46.055 49.65 46.265 ;
		RECT	49.11 46.38 49.65 46.57 ;
		RECT	49.11 47.245 49.65 47.435 ;
		RECT	49.11 48.03 49.65 48.13 ;
		RECT	49.11 48.52 49.65 48.62 ;
		RECT	49.11 49.01 49.65 49.115 ;
		RECT	49.11 49.505 49.65 49.605 ;
		RECT	49.11 49.995 49.65 50.1 ;
		RECT	49.11 50.69 49.65 50.88 ;
		RECT	49.11 51.495 49.65 51.685 ;
		RECT	49.11 51.83 49.65 52.04 ;
		RECT	49.11 52.47 49.65 52.555 ;
		RECT	49.11 52.945 49.65 53.05 ;
		RECT	49.11 53.44 49.65 53.545 ;
		RECT	49.11 53.935 49.65 54.025 ;
		RECT	49.11 54.435 49.65 54.515 ;
		RECT	49.11 54.615 49.65 54.825 ;
		RECT	49.11 54.925 49.65 55.02 ;
		RECT	49.11 55.41 49.65 55.51 ;
		RECT	49.11 55.9 49.65 56.005 ;
		RECT	49.11 56.395 49.65 56.485 ;
		RECT	49.11 56.895 49.65 56.985 ;
		RECT	49.11 57.375 49.65 57.48 ;
		RECT	49.11 57.87 49.65 57.97 ;
		RECT	49.11 58.36 49.65 58.465 ;
		RECT	49.11 58.565 49.65 58.755 ;
		RECT	49.11 58.855 49.65 58.955 ;
		RECT	49.11 59.345 49.65 59.445 ;
		RECT	49.11 59.835 49.65 59.94 ;
		RECT	49.11 60.33 49.65 60.43 ;
		RECT	49.11 60.82 49.65 60.925 ;
		RECT	49.11 61.315 49.65 61.415 ;
		RECT	49.11 61.805 49.65 61.905 ;
		RECT	49.11 62.49 49.65 62.7 ;
		RECT	49.11 62.8 49.65 62.89 ;
		RECT	49.11 63.28 49.65 63.375 ;
		RECT	49.11 63.79 49.65 63.86 ;
		RECT	49.11 64.28 49.65 64.35 ;
		RECT	49.11 64.765 49.65 64.825 ;
		RECT	49.11 65.215 49.65 65.35 ;
		RECT	49.11 65.74 49.65 65.81 ;
		RECT	49.11 66.2 49.65 66.35 ;
		RECT	49.11 66.45 49.65 66.64 ;
		RECT	49.11 66.925 49.65 67.115 ;
		RECT	49.11 67.215 49.65 67.32 ;
		RECT	49.11 68.2 49.65 68.305 ;
		RECT	49.11 68.705 49.65 68.915 ;
		RECT	49.65 29.15 50.25 29.34 ;
		RECT	49.65 29.825 50.25 29.925 ;
		RECT	49.65 30.805 50.25 30.91 ;
		RECT	49.65 31.01 50.25 31.2 ;
		RECT	49.65 31.485 50.25 31.675 ;
		RECT	49.65 31.78 50.415 31.93 ;
		RECT	49.65 32.32 50.25 32.385 ;
		RECT	49.65 32.775 50.25 32.88 ;
		RECT	49.65 33.27 50.25 33.37 ;
		RECT	49.65 34.25 50.25 34.355 ;
		RECT	49.65 34.745 50.25 34.845 ;
		RECT	49.65 35.235 50.25 35.34 ;
		RECT	49.65 35.44 50.25 35.63 ;
		RECT	49.65 35.73 50.25 35.83 ;
		RECT	49.65 36.22 50.25 36.325 ;
		RECT	49.65 36.715 50.25 36.815 ;
		RECT	49.65 37.205 50.25 37.305 ;
		RECT	49.65 37.695 50.25 37.8 ;
		RECT	49.65 38.19 50.25 38.29 ;
		RECT	49.65 38.68 50.25 38.78 ;
		RECT	49.65 39.17 50.25 39.275 ;
		RECT	49.65 39.375 50.25 39.565 ;
		RECT	49.65 39.665 50.25 39.765 ;
		RECT	49.65 40.155 50.25 40.26 ;
		RECT	49.65 40.65 50.25 40.75 ;
		RECT	49.65 41.14 50.25 41.23 ;
		RECT	49.65 41.64 50.25 41.735 ;
		RECT	49.65 42.125 50.25 42.225 ;
		RECT	49.65 42.615 50.25 42.72 ;
		RECT	49.65 43.11 50.25 43.2 ;
		RECT	49.65 43.3 50.25 43.51 ;
		RECT	49.65 43.61 50.25 43.705 ;
		RECT	49.65 44.095 50.25 44.2 ;
		RECT	49.65 44.59 50.25 44.685 ;
		RECT	49.65 45.075 50.25 45.18 ;
		RECT	49.65 45.57 50.25 45.655 ;
		RECT	49.65 46.055 50.325 46.265 ;
		RECT	49.65 46.38 50.25 46.57 ;
		RECT	49.65 47.245 50.25 47.435 ;
		RECT	49.65 48.03 50.25 48.13 ;
		RECT	49.65 48.52 50.25 48.62 ;
		RECT	49.65 49.01 50.25 49.115 ;
		RECT	49.65 49.505 50.25 49.605 ;
		RECT	49.65 49.995 50.25 50.1 ;
		RECT	49.65 50.69 50.25 50.88 ;
		RECT	49.65 51.495 50.25 51.685 ;
		RECT	49.65 51.83 50.25 52.04 ;
		RECT	49.65 52.47 50.25 52.555 ;
		RECT	49.65 52.945 50.25 53.05 ;
		RECT	49.65 53.44 50.25 53.545 ;
		RECT	49.65 53.935 50.25 54.025 ;
		RECT	49.65 54.435 50.25 54.515 ;
		RECT	49.65 54.615 50.25 54.825 ;
		RECT	49.65 54.925 50.25 55.02 ;
		RECT	49.65 55.41 50.25 55.51 ;
		RECT	49.65 55.9 50.25 56.005 ;
		RECT	49.65 56.395 50.25 56.485 ;
		RECT	49.65 56.895 50.25 56.985 ;
		RECT	49.65 57.375 50.25 57.48 ;
		RECT	49.65 57.87 50.25 57.97 ;
		RECT	49.65 58.36 50.25 58.465 ;
		RECT	49.65 58.565 50.25 58.755 ;
		RECT	49.65 58.855 50.25 58.955 ;
		RECT	49.65 59.345 50.25 59.445 ;
		RECT	49.65 59.835 50.25 59.94 ;
		RECT	49.65 60.33 50.25 60.43 ;
		RECT	49.65 60.82 50.25 60.925 ;
		RECT	49.65 61.315 50.25 61.415 ;
		RECT	49.65 61.805 50.25 61.905 ;
		RECT	49.65 62.49 50.25 62.7 ;
		RECT	49.65 62.8 50.25 62.89 ;
		RECT	49.65 63.28 50.25 63.375 ;
		RECT	49.65 63.79 50.25 63.86 ;
		RECT	49.65 64.28 50.25 64.35 ;
		RECT	49.65 64.765 50.25 64.825 ;
		RECT	49.65 65.215 50.25 65.35 ;
		RECT	49.65 65.74 50.25 65.81 ;
		RECT	49.65 66.2 50.25 66.35 ;
		RECT	49.65 66.45 50.25 66.64 ;
		RECT	49.65 66.925 50.25 67.115 ;
		RECT	49.65 67.215 50.25 67.32 ;
		RECT	49.65 68.2 50.25 68.305 ;
		RECT	49.65 68.705 50.25 68.915 ;
		RECT	0.295 34.455 50.93 34.645 ;
		RECT	0.215 43.805 51.11 43.995 ;
		RECT	0.21 45.755 51.1 45.945 ;
		RECT	0.22 52.18 51.11 52.37 ;
		RECT	0.225 54.125 51.11 54.335 ;
		RECT	0.225 63.475 50.93 63.685 ;
		RECT	0.225 63.79 0.57 63.86 ;
		RECT	0.22 64.28 0.57 64.35 ;
		RECT	11.61 30.32 51.31 30.41 ;
		RECT	11.61 31.305 51.31 31.385 ;
		RECT	14.2 33.765 50.6 33.855 ;
		RECT	13.85 47.05 51.31 47.14 ;
		RECT	13.85 47.545 51.31 47.635 ;
		RECT	7.07 49.015 13.545 49.115 ;
		RECT	13.85 50.495 51.31 50.585 ;
		RECT	13.85 50.985 51.31 51.075 ;
		RECT	14.2 62.3 50.6 62.39 ;
		RECT	0.57 62.805 2.735 62.875 ;
		RECT	12.605 66.74 51.31 66.82 ;
		RECT	12.605 67.715 51.31 67.805 ;
		RECT	50.25 63.79 50.93 63.86 ;
		RECT	50.25 64.28 50.93 64.35 ;
		LAYER	VIA1 DESIGNRULEWIDTH 0.07 ;
		RECT	0 0 51.405 100.94 ;
		LAYER	VIA2 DESIGNRULEWIDTH 0.07 ;
		RECT	0 0 51.405 100.94 ;
		LAYER	VIA3 DESIGNRULEWIDTH 0.07 ;
		RECT	0.435 28.015 0.485 28.145 ;
		RECT	0.435 29.18 0.485 29.31 ;
		RECT	0.435 31.045 0.485 31.175 ;
		RECT	0.435 31.515 0.485 31.645 ;
		RECT	0.435 35.47 0.485 35.6 ;
		RECT	0.435 39.405 0.485 39.535 ;
		RECT	0.435 43.34 0.485 43.47 ;
		RECT	0.435 46.465 0.485 46.595 ;
		RECT	0.435 47.275 0.485 47.405 ;
		RECT	0.435 50.72 0.485 50.85 ;
		RECT	0.435 51.53 0.485 51.66 ;
		RECT	0.435 54.655 0.485 54.785 ;
		RECT	0.435 58.595 0.485 58.725 ;
		RECT	0.435 62.53 0.485 62.66 ;
		RECT	0.435 66.48 0.485 66.61 ;
		RECT	0.435 66.955 0.485 67.085 ;
		RECT	0.435 68.745 0.485 68.875 ;
		RECT	0.435 69.915 0.485 70.045 ;
		RECT	0.435 28.475 0.485 28.605 ;
		RECT	0.435 34.485 0.485 34.615 ;
		RECT	0.435 63.515 0.485 63.645 ;
		RECT	0.435 69.455 0.485 69.585 ;
		RECT	1.085 28.015 1.135 28.145 ;
		RECT	1.38 28.015 1.43 28.145 ;
		RECT	1.86 28.015 1.91 28.145 ;
		RECT	2.01 28.015 2.06 28.145 ;
		RECT	3.25 28.015 3.3 28.145 ;
		RECT	3.515 28.015 3.565 28.145 ;
		RECT	4.51 28.015 4.56 28.145 ;
		RECT	5.035 28.015 5.085 28.145 ;
		RECT	6.22 28.015 6.27 28.145 ;
		RECT	7.5 28.015 7.55 28.145 ;
		RECT	9.315 28.015 9.365 28.145 ;
		RECT	9.72 28.015 9.77 28.145 ;
		RECT	11.025 28.015 11.075 28.145 ;
		RECT	0.62 28.245 0.67 28.375 ;
		RECT	3.65 28.245 3.7 28.375 ;
		RECT	7.19 28.245 7.24 28.375 ;
		RECT	14.14 28.245 14.19 28.375 ;
		RECT	2.18 28.475 2.23 28.605 ;
		RECT	8.56 28.475 8.61 28.605 ;
		RECT	10.27 28.475 10.32 28.605 ;
		RECT	13.8 28.705 13.85 28.835 ;
		RECT	1.045 29.155 1.175 29.205 ;
		RECT	1.34 29.155 1.47 29.205 ;
		RECT	4.47 29.155 4.6 29.205 ;
		RECT	9.275 29.155 9.405 29.205 ;
		RECT	1.86 29.18 1.91 29.31 ;
		RECT	2.01 29.18 2.06 29.31 ;
		RECT	3.25 29.18 3.3 29.31 ;
		RECT	3.515 29.18 3.565 29.31 ;
		RECT	5.035 29.18 5.085 29.31 ;
		RECT	6.22 29.18 6.27 29.31 ;
		RECT	7.5 29.18 7.55 29.31 ;
		RECT	9.72 29.18 9.77 29.31 ;
		RECT	11.025 29.18 11.075 29.31 ;
		RECT	1.045 29.285 1.175 29.335 ;
		RECT	1.34 29.285 1.47 29.335 ;
		RECT	4.47 29.285 4.6 29.335 ;
		RECT	9.275 29.285 9.405 29.335 ;
		RECT	3.02 29.54 3.15 29.59 ;
		RECT	1.57 29.565 1.62 29.695 ;
		RECT	4.87 29.565 4.92 29.695 ;
		RECT	5.9 29.565 5.95 29.695 ;
		RECT	8.955 29.565 9.005 29.695 ;
		RECT	12.79 29.565 12.84 29.695 ;
		RECT	14.33 29.565 14.38 29.695 ;
		RECT	3.02 29.67 3.15 29.72 ;
		RECT	3.8 30.03 3.93 30.08 ;
		RECT	5.635 30.03 5.765 30.08 ;
		RECT	8.31 30.03 8.44 30.08 ;
		RECT	8.73 30.03 8.86 30.08 ;
		RECT	0.9 30.055 0.95 30.185 ;
		RECT	2.485 30.055 2.535 30.185 ;
		RECT	2.615 30.055 2.665 30.185 ;
		RECT	6.065 30.055 6.115 30.185 ;
		RECT	6.725 30.055 6.775 30.185 ;
		RECT	11.555 30.055 11.865 30.185 ;
		RECT	12.52 30.055 12.57 30.185 ;
		RECT	14.005 30.055 14.055 30.185 ;
		RECT	3.8 30.16 3.93 30.21 ;
		RECT	5.635 30.16 5.765 30.21 ;
		RECT	8.31 30.16 8.44 30.21 ;
		RECT	8.73 30.16 8.86 30.21 ;
		RECT	11.685 30.34 11.735 30.39 ;
		RECT	12.655 30.34 12.705 30.39 ;
		RECT	3.02 30.52 3.15 30.57 ;
		RECT	1.57 30.545 1.62 30.675 ;
		RECT	4.87 30.545 4.92 30.675 ;
		RECT	5.9 30.545 5.95 30.675 ;
		RECT	8.955 30.545 9.005 30.675 ;
		RECT	12.79 30.545 12.84 30.675 ;
		RECT	14.335 30.545 14.385 30.675 ;
		RECT	3.02 30.65 3.15 30.7 ;
		RECT	1.045 31.02 1.175 31.07 ;
		RECT	1.34 31.02 1.47 31.07 ;
		RECT	4.47 31.02 4.6 31.07 ;
		RECT	9.275 31.02 9.405 31.07 ;
		RECT	13.675 31.04 13.725 31.17 ;
		RECT	1.86 31.045 1.91 31.175 ;
		RECT	2.01 31.045 2.06 31.175 ;
		RECT	3.25 31.045 3.3 31.175 ;
		RECT	3.515 31.045 3.565 31.175 ;
		RECT	5.035 31.045 5.085 31.175 ;
		RECT	6.22 31.045 6.27 31.175 ;
		RECT	7.5 31.045 7.55 31.175 ;
		RECT	9.72 31.045 9.77 31.175 ;
		RECT	11.025 31.045 11.075 31.175 ;
		RECT	1.045 31.15 1.175 31.2 ;
		RECT	1.34 31.15 1.47 31.2 ;
		RECT	4.47 31.15 4.6 31.2 ;
		RECT	9.275 31.15 9.405 31.2 ;
		RECT	11.685 31.32 11.735 31.37 ;
		RECT	12.655 31.32 12.705 31.37 ;
		RECT	1.045 31.49 1.175 31.54 ;
		RECT	1.34 31.49 1.47 31.54 ;
		RECT	4.47 31.49 4.6 31.54 ;
		RECT	9.275 31.49 9.405 31.54 ;
		RECT	1.86 31.515 1.91 31.645 ;
		RECT	2.01 31.515 2.06 31.645 ;
		RECT	3.25 31.515 3.3 31.645 ;
		RECT	3.515 31.515 3.565 31.645 ;
		RECT	5.035 31.515 5.085 31.645 ;
		RECT	6.22 31.515 6.27 31.645 ;
		RECT	7.5 31.515 7.55 31.645 ;
		RECT	9.72 31.515 9.77 31.645 ;
		RECT	11.025 31.515 11.075 31.645 ;
		RECT	1.045 31.62 1.175 31.67 ;
		RECT	1.34 31.62 1.47 31.67 ;
		RECT	4.47 31.62 4.6 31.67 ;
		RECT	9.275 31.62 9.405 31.67 ;
		RECT	3.8 32.035 3.93 32.085 ;
		RECT	5.635 32.035 5.765 32.085 ;
		RECT	8.31 32.035 8.44 32.085 ;
		RECT	8.73 32.035 8.86 32.085 ;
		RECT	0.9 32.06 0.95 32.19 ;
		RECT	2.485 32.06 2.535 32.19 ;
		RECT	2.615 32.06 2.665 32.19 ;
		RECT	6.065 32.06 6.115 32.19 ;
		RECT	6.725 32.06 6.775 32.19 ;
		RECT	11.555 32.06 11.865 32.19 ;
		RECT	12.52 32.06 12.57 32.19 ;
		RECT	14.005 32.06 14.055 32.19 ;
		RECT	3.8 32.165 3.93 32.215 ;
		RECT	5.635 32.165 5.765 32.215 ;
		RECT	8.31 32.165 8.44 32.215 ;
		RECT	8.73 32.165 8.86 32.215 ;
		RECT	3.02 32.49 3.15 32.54 ;
		RECT	1.57 32.515 1.62 32.645 ;
		RECT	4.87 32.515 4.92 32.645 ;
		RECT	5.9 32.515 5.95 32.645 ;
		RECT	8.955 32.515 9.005 32.645 ;
		RECT	12.79 32.515 12.84 32.645 ;
		RECT	14.335 32.515 14.385 32.645 ;
		RECT	3.02 32.62 3.15 32.67 ;
		RECT	4.035 33.01 4.085 33.14 ;
		RECT	6.495 33.01 6.545 33.14 ;
		RECT	11.685 33.01 11.735 33.14 ;
		RECT	12.655 33.01 12.705 33.14 ;
		RECT	3.02 33.475 3.15 33.525 ;
		RECT	1.57 33.5 1.62 33.63 ;
		RECT	4.87 33.5 4.92 33.63 ;
		RECT	5.9 33.5 5.95 33.63 ;
		RECT	8.955 33.5 9.005 33.63 ;
		RECT	12.79 33.5 12.84 33.63 ;
		RECT	14.335 33.5 14.385 33.63 ;
		RECT	3.02 33.605 3.15 33.655 ;
		RECT	14.29 33.785 14.42 33.835 ;
		RECT	4.035 33.99 4.085 34.12 ;
		RECT	6.495 33.99 6.545 34.12 ;
		RECT	2.18 34.485 2.23 34.615 ;
		RECT	8.56 34.485 8.61 34.615 ;
		RECT	10.27 34.485 10.32 34.615 ;
		RECT	3.8 34.95 3.93 35 ;
		RECT	5.635 34.95 5.765 35 ;
		RECT	8.31 34.95 8.44 35 ;
		RECT	8.73 34.95 8.86 35 ;
		RECT	0.9 34.975 0.95 35.105 ;
		RECT	2.485 34.975 2.535 35.105 ;
		RECT	2.615 34.975 2.665 35.105 ;
		RECT	6.065 34.975 6.115 35.105 ;
		RECT	6.725 34.975 6.775 35.105 ;
		RECT	11.555 34.975 11.865 35.105 ;
		RECT	12.52 34.975 12.57 35.105 ;
		RECT	14.005 34.975 14.055 35.105 ;
		RECT	3.8 35.08 3.93 35.13 ;
		RECT	5.635 35.08 5.765 35.13 ;
		RECT	8.31 35.08 8.44 35.13 ;
		RECT	8.73 35.08 8.86 35.13 ;
		RECT	1.045 35.445 1.175 35.495 ;
		RECT	1.34 35.445 1.47 35.495 ;
		RECT	4.47 35.445 4.6 35.495 ;
		RECT	1.86 35.47 1.91 35.6 ;
		RECT	2.01 35.47 2.06 35.6 ;
		RECT	2.32 35.47 2.37 35.6 ;
		RECT	3.25 35.47 3.3 35.6 ;
		RECT	3.515 35.47 3.565 35.6 ;
		RECT	5.035 35.47 5.085 35.6 ;
		RECT	6.22 35.47 6.27 35.6 ;
		RECT	7.5 35.47 7.55 35.6 ;
		RECT	9.72 35.47 9.77 35.6 ;
		RECT	11.025 35.47 11.075 35.6 ;
		RECT	1.045 35.575 1.175 35.625 ;
		RECT	1.34 35.575 1.47 35.625 ;
		RECT	4.47 35.575 4.6 35.625 ;
		RECT	3.8 35.935 3.93 35.985 ;
		RECT	5.635 35.935 5.765 35.985 ;
		RECT	8.31 35.935 8.44 35.985 ;
		RECT	8.73 35.935 8.86 35.985 ;
		RECT	0.9 35.96 0.95 36.09 ;
		RECT	2.485 35.96 2.535 36.09 ;
		RECT	2.615 35.96 2.665 36.09 ;
		RECT	6.065 35.96 6.115 36.09 ;
		RECT	6.725 35.96 6.775 36.09 ;
		RECT	11.555 35.96 11.865 36.09 ;
		RECT	12.52 35.96 12.57 36.09 ;
		RECT	14.005 35.96 14.055 36.09 ;
		RECT	3.8 36.065 3.93 36.115 ;
		RECT	5.635 36.065 5.765 36.115 ;
		RECT	8.31 36.065 8.44 36.115 ;
		RECT	8.73 36.065 8.86 36.115 ;
		RECT	3.02 36.43 3.15 36.48 ;
		RECT	1.57 36.455 1.62 36.585 ;
		RECT	4.87 36.455 4.92 36.585 ;
		RECT	5.9 36.455 5.95 36.585 ;
		RECT	9.195 36.455 9.245 36.585 ;
		RECT	10.27 36.455 10.32 36.585 ;
		RECT	12.79 36.455 12.84 36.585 ;
		RECT	14.335 36.455 14.385 36.585 ;
		RECT	3.02 36.56 3.15 36.61 ;
		RECT	4.035 36.945 4.085 37.075 ;
		RECT	3.02 37.41 3.15 37.46 ;
		RECT	1.57 37.435 1.62 37.565 ;
		RECT	4.87 37.435 4.92 37.565 ;
		RECT	5.9 37.435 5.95 37.565 ;
		RECT	9.195 37.435 9.245 37.565 ;
		RECT	9.43 37.435 9.48 37.565 ;
		RECT	10.27 37.435 10.32 37.565 ;
		RECT	12.79 37.435 12.84 37.565 ;
		RECT	14.335 37.435 14.385 37.565 ;
		RECT	3.02 37.54 3.15 37.59 ;
		RECT	0.9 37.905 14.055 38.085 ;
		RECT	3.02 38.395 3.15 38.445 ;
		RECT	1.57 38.42 1.62 38.55 ;
		RECT	4.87 38.42 4.92 38.55 ;
		RECT	5.9 38.42 5.95 38.55 ;
		RECT	9.43 38.42 9.48 38.55 ;
		RECT	10.27 38.42 10.32 38.55 ;
		RECT	12.79 38.42 12.84 38.55 ;
		RECT	14.33 38.42 14.38 38.55 ;
		RECT	3.02 38.525 3.15 38.575 ;
		RECT	3.8 38.885 3.93 38.935 ;
		RECT	5.635 38.885 5.765 38.935 ;
		RECT	8.31 38.885 8.44 38.935 ;
		RECT	8.73 38.885 8.86 38.935 ;
		RECT	0.9 38.91 0.95 39.04 ;
		RECT	2.485 38.91 2.535 39.04 ;
		RECT	2.615 38.91 2.665 39.04 ;
		RECT	6.065 38.91 6.115 39.04 ;
		RECT	6.725 38.91 6.775 39.04 ;
		RECT	11.555 38.91 11.865 39.04 ;
		RECT	12.52 38.91 12.57 39.04 ;
		RECT	14.005 38.91 14.055 39.04 ;
		RECT	3.8 39.015 3.93 39.065 ;
		RECT	5.635 39.015 5.765 39.065 ;
		RECT	8.31 39.015 8.44 39.065 ;
		RECT	8.73 39.015 8.86 39.065 ;
		RECT	1.045 39.38 1.175 39.43 ;
		RECT	1.34 39.38 1.47 39.43 ;
		RECT	4.47 39.38 4.6 39.43 ;
		RECT	1.86 39.405 1.91 39.535 ;
		RECT	2.01 39.405 2.06 39.535 ;
		RECT	2.32 39.405 2.37 39.535 ;
		RECT	3.25 39.405 3.3 39.535 ;
		RECT	3.515 39.405 3.565 39.535 ;
		RECT	5.035 39.405 5.085 39.535 ;
		RECT	6.22 39.405 6.27 39.535 ;
		RECT	7.5 39.405 7.55 39.535 ;
		RECT	9.72 39.405 9.77 39.535 ;
		RECT	11.025 39.405 11.075 39.535 ;
		RECT	1.045 39.51 1.175 39.56 ;
		RECT	1.34 39.51 1.47 39.56 ;
		RECT	4.47 39.51 4.6 39.56 ;
		RECT	3.8 39.87 3.93 39.92 ;
		RECT	5.635 39.87 5.765 39.92 ;
		RECT	8.31 39.87 8.44 39.92 ;
		RECT	8.73 39.87 8.86 39.92 ;
		RECT	0.9 39.895 0.95 40.025 ;
		RECT	2.485 39.895 2.535 40.025 ;
		RECT	2.615 39.895 2.665 40.025 ;
		RECT	6.065 39.895 6.115 40.025 ;
		RECT	6.725 39.895 6.775 40.025 ;
		RECT	11.555 39.895 11.865 40.025 ;
		RECT	12.52 39.895 12.57 40.025 ;
		RECT	14.005 39.895 14.055 40.025 ;
		RECT	3.8 40 3.93 40.05 ;
		RECT	5.635 40 5.765 40.05 ;
		RECT	8.31 40 8.44 40.05 ;
		RECT	8.73 40 8.86 40.05 ;
		RECT	3.02 40.365 3.15 40.415 ;
		RECT	1.57 40.39 1.62 40.52 ;
		RECT	4.87 40.39 4.92 40.52 ;
		RECT	5.9 40.39 5.95 40.52 ;
		RECT	6.375 40.39 6.425 40.52 ;
		RECT	10.27 40.39 10.32 40.52 ;
		RECT	12.65 40.39 12.84 40.52 ;
		RECT	14.33 40.39 14.38 40.52 ;
		RECT	3.02 40.495 3.15 40.545 ;
		RECT	4.035 40.88 4.085 41.01 ;
		RECT	6.835 41.165 6.885 41.215 ;
		RECT	3.02 41.345 3.15 41.395 ;
		RECT	1.57 41.37 1.62 41.5 ;
		RECT	4.87 41.37 4.92 41.5 ;
		RECT	5.9 41.37 5.95 41.5 ;
		RECT	6.375 41.37 6.425 41.5 ;
		RECT	7.015 41.37 7.065 41.5 ;
		RECT	10.27 41.37 10.32 41.5 ;
		RECT	12.79 41.37 12.84 41.5 ;
		RECT	14.33 41.37 14.38 41.5 ;
		RECT	3.02 41.475 3.15 41.525 ;
		RECT	4.035 41.865 4.085 41.995 ;
		RECT	3.02 42.33 3.15 42.38 ;
		RECT	1.57 42.355 1.62 42.485 ;
		RECT	4.87 42.355 4.92 42.485 ;
		RECT	5.9 42.355 5.95 42.485 ;
		RECT	6.375 42.355 6.425 42.485 ;
		RECT	7.015 42.355 7.065 42.485 ;
		RECT	10.27 42.355 10.32 42.485 ;
		RECT	12.79 42.355 12.84 42.485 ;
		RECT	14.33 42.355 14.38 42.485 ;
		RECT	3.02 42.46 3.15 42.51 ;
		RECT	0.9 42.85 0.95 42.98 ;
		RECT	2.485 42.85 2.535 42.98 ;
		RECT	2.615 42.85 2.665 42.98 ;
		RECT	6.065 42.85 6.115 42.98 ;
		RECT	6.675 42.85 6.725 42.98 ;
		RECT	11.555 42.85 11.865 42.98 ;
		RECT	12.52 42.85 12.57 42.98 ;
		RECT	14.005 42.85 14.055 42.98 ;
		RECT	3.8 42.89 3.93 42.94 ;
		RECT	5.635 42.89 5.765 42.94 ;
		RECT	8.31 42.89 8.44 42.94 ;
		RECT	8.73 42.89 8.86 42.94 ;
		RECT	9.315 43.135 9.445 43.185 ;
		RECT	1.045 43.315 1.175 43.365 ;
		RECT	1.34 43.315 1.47 43.365 ;
		RECT	4.47 43.315 4.6 43.365 ;
		RECT	1.86 43.34 1.91 43.47 ;
		RECT	2.01 43.34 2.06 43.47 ;
		RECT	2.32 43.34 2.37 43.47 ;
		RECT	3.25 43.34 3.3 43.47 ;
		RECT	3.515 43.34 3.565 43.47 ;
		RECT	5.035 43.34 5.085 43.47 ;
		RECT	6.22 43.34 6.27 43.47 ;
		RECT	7.5 43.34 7.55 43.47 ;
		RECT	9.72 43.34 9.77 43.47 ;
		RECT	11.025 43.34 11.075 43.47 ;
		RECT	1.045 43.445 1.175 43.495 ;
		RECT	1.34 43.445 1.47 43.495 ;
		RECT	4.47 43.445 4.6 43.495 ;
		RECT	0.62 43.835 0.67 43.965 ;
		RECT	3.65 43.835 3.7 43.965 ;
		RECT	7.19 43.835 7.24 43.965 ;
		RECT	14.14 43.835 14.19 43.965 ;
		RECT	3.02 44.305 3.15 44.355 ;
		RECT	1.57 44.33 1.62 44.46 ;
		RECT	4.87 44.33 4.92 44.46 ;
		RECT	5.9 44.33 5.95 44.46 ;
		RECT	6.375 44.33 6.425 44.46 ;
		RECT	7.015 44.33 7.065 44.46 ;
		RECT	10.27 44.33 10.32 44.46 ;
		RECT	12.79 44.33 12.84 44.46 ;
		RECT	14.335 44.33 14.385 44.46 ;
		RECT	3.02 44.435 3.15 44.485 ;
		RECT	4.035 44.815 4.085 44.945 ;
		RECT	11.685 44.815 11.735 44.945 ;
		RECT	13.9 44.815 13.95 44.945 ;
		RECT	3.02 45.285 3.15 45.335 ;
		RECT	1.57 45.31 1.62 45.44 ;
		RECT	4.87 45.31 4.92 45.44 ;
		RECT	5.9 45.31 5.95 45.44 ;
		RECT	6.375 45.31 6.425 45.44 ;
		RECT	7.015 45.31 7.065 45.44 ;
		RECT	10.27 45.31 10.32 45.44 ;
		RECT	12.79 45.31 12.84 45.44 ;
		RECT	14.335 45.31 14.385 45.44 ;
		RECT	3.02 45.415 3.15 45.465 ;
		RECT	13.8 45.785 13.85 45.915 ;
		RECT	13.675 46.41 13.725 46.54 ;
		RECT	1.085 46.465 1.135 46.595 ;
		RECT	1.38 46.465 1.43 46.595 ;
		RECT	1.86 46.465 1.91 46.595 ;
		RECT	2.01 46.465 2.06 46.595 ;
		RECT	2.32 46.465 2.37 46.595 ;
		RECT	3.25 46.465 3.3 46.595 ;
		RECT	3.515 46.465 3.565 46.595 ;
		RECT	4.51 46.465 4.56 46.595 ;
		RECT	5.035 46.465 5.085 46.595 ;
		RECT	6.22 46.465 6.27 46.595 ;
		RECT	7.5 46.465 7.55 46.595 ;
		RECT	9.72 46.465 9.77 46.595 ;
		RECT	11.025 46.465 11.075 46.595 ;
		RECT	3.8 46.76 3.93 46.81 ;
		RECT	5.635 46.76 5.765 46.81 ;
		RECT	8.31 46.76 8.44 46.81 ;
		RECT	8.73 46.76 8.86 46.81 ;
		RECT	0.9 46.785 0.95 46.915 ;
		RECT	2.485 46.785 2.535 46.915 ;
		RECT	2.615 46.785 2.665 46.915 ;
		RECT	6.065 46.785 6.115 46.915 ;
		RECT	6.675 46.785 6.725 46.915 ;
		RECT	11.555 46.785 11.865 46.915 ;
		RECT	12.52 46.785 12.57 46.915 ;
		RECT	14.005 46.785 14.055 46.915 ;
		RECT	3.8 46.89 3.93 46.94 ;
		RECT	5.635 46.89 5.765 46.94 ;
		RECT	8.31 46.89 8.44 46.94 ;
		RECT	8.73 46.89 8.86 46.94 ;
		RECT	13.9 47.07 13.95 47.12 ;
		RECT	1.045 47.25 1.175 47.3 ;
		RECT	1.34 47.25 1.47 47.3 ;
		RECT	4.47 47.25 4.6 47.3 ;
		RECT	1.86 47.275 1.91 47.405 ;
		RECT	2.01 47.275 2.06 47.405 ;
		RECT	2.32 47.275 2.37 47.405 ;
		RECT	3.25 47.275 3.3 47.405 ;
		RECT	3.515 47.275 3.565 47.405 ;
		RECT	5.035 47.275 5.085 47.405 ;
		RECT	6.22 47.275 6.27 47.405 ;
		RECT	7.5 47.275 7.55 47.405 ;
		RECT	9.72 47.275 9.77 47.405 ;
		RECT	11.025 47.275 11.075 47.405 ;
		RECT	1.045 47.38 1.175 47.43 ;
		RECT	1.34 47.38 1.47 47.43 ;
		RECT	4.47 47.38 4.6 47.43 ;
		RECT	13.9 47.565 13.95 47.615 ;
		RECT	3.8 47.745 3.93 47.795 ;
		RECT	5.635 47.745 5.765 47.795 ;
		RECT	8.31 47.745 8.44 47.795 ;
		RECT	8.73 47.745 8.86 47.795 ;
		RECT	0.9 47.77 0.95 47.9 ;
		RECT	2.485 47.77 2.535 47.9 ;
		RECT	2.615 47.77 2.665 47.9 ;
		RECT	6.065 47.77 6.115 47.9 ;
		RECT	6.675 47.77 6.725 47.9 ;
		RECT	10.12 47.77 10.17 47.9 ;
		RECT	11.555 47.77 11.865 47.9 ;
		RECT	12.52 47.77 12.57 47.9 ;
		RECT	14.005 47.77 14.055 47.9 ;
		RECT	3.8 47.875 3.93 47.925 ;
		RECT	5.635 47.875 5.765 47.925 ;
		RECT	8.31 47.875 8.44 47.925 ;
		RECT	8.73 47.875 8.86 47.925 ;
		RECT	3.02 48.235 3.15 48.285 ;
		RECT	1.57 48.26 1.62 48.39 ;
		RECT	4.87 48.26 4.92 48.39 ;
		RECT	5.9 48.26 5.95 48.39 ;
		RECT	6.375 48.26 6.425 48.39 ;
		RECT	7.015 48.26 7.065 48.39 ;
		RECT	9.11 48.26 9.16 48.39 ;
		RECT	10.27 48.26 10.32 48.39 ;
		RECT	12.79 48.26 12.84 48.39 ;
		RECT	14.335 48.26 14.385 48.39 ;
		RECT	3.02 48.365 3.15 48.415 ;
		RECT	4.035 48.75 4.085 48.88 ;
		RECT	13.9 48.75 13.95 48.88 ;
		RECT	7.19 49.04 7.24 49.09 ;
		RECT	12.655 49.04 12.705 49.09 ;
		RECT	4.035 49.245 4.085 49.375 ;
		RECT	13.9 49.245 13.95 49.375 ;
		RECT	3.02 49.71 3.15 49.76 ;
		RECT	1.57 49.735 1.62 49.865 ;
		RECT	4.87 49.735 4.92 49.865 ;
		RECT	5.9 49.735 5.95 49.865 ;
		RECT	6.375 49.735 6.425 49.865 ;
		RECT	7.015 49.735 7.065 49.865 ;
		RECT	9.11 49.735 9.16 49.865 ;
		RECT	10.27 49.735 10.32 49.865 ;
		RECT	12.79 49.735 12.84 49.865 ;
		RECT	14.335 49.735 14.385 49.865 ;
		RECT	3.02 49.84 3.15 49.89 ;
		RECT	3.8 50.205 3.93 50.255 ;
		RECT	4.22 50.205 4.35 50.255 ;
		RECT	5.635 50.205 5.765 50.255 ;
		RECT	8.31 50.205 8.44 50.255 ;
		RECT	8.73 50.205 8.86 50.255 ;
		RECT	0.9 50.23 0.95 50.36 ;
		RECT	2.485 50.23 2.535 50.36 ;
		RECT	2.615 50.23 2.665 50.36 ;
		RECT	6.065 50.23 6.115 50.36 ;
		RECT	6.675 50.23 6.725 50.36 ;
		RECT	10.12 50.23 10.17 50.36 ;
		RECT	11.555 50.23 11.865 50.36 ;
		RECT	12.52 50.23 12.57 50.36 ;
		RECT	14.005 50.23 14.055 50.36 ;
		RECT	3.8 50.335 3.93 50.385 ;
		RECT	4.22 50.335 4.35 50.385 ;
		RECT	5.635 50.335 5.765 50.385 ;
		RECT	8.31 50.335 8.44 50.385 ;
		RECT	8.73 50.335 8.86 50.385 ;
		RECT	13.9 50.515 13.95 50.565 ;
		RECT	1.045 50.695 1.175 50.745 ;
		RECT	1.34 50.695 1.47 50.745 ;
		RECT	4.47 50.695 4.6 50.745 ;
		RECT	1.86 50.72 1.91 50.85 ;
		RECT	2.01 50.72 2.06 50.85 ;
		RECT	2.32 50.72 2.37 50.85 ;
		RECT	3.25 50.72 3.3 50.85 ;
		RECT	3.515 50.72 3.565 50.85 ;
		RECT	5.035 50.72 5.085 50.85 ;
		RECT	6.22 50.72 6.27 50.85 ;
		RECT	7.5 50.72 7.55 50.85 ;
		RECT	9.72 50.72 9.77 50.85 ;
		RECT	11.025 50.72 11.075 50.85 ;
		RECT	1.045 50.825 1.175 50.875 ;
		RECT	1.34 50.825 1.47 50.875 ;
		RECT	4.47 50.825 4.6 50.875 ;
		RECT	13.9 51.005 13.95 51.055 ;
		RECT	0.9 51.185 14.055 51.365 ;
		RECT	13.675 51.525 13.725 51.655 ;
		RECT	1.085 51.53 1.135 51.66 ;
		RECT	1.38 51.53 1.43 51.66 ;
		RECT	1.86 51.53 1.91 51.66 ;
		RECT	2.01 51.53 2.06 51.66 ;
		RECT	2.32 51.53 2.37 51.66 ;
		RECT	3.25 51.53 3.3 51.66 ;
		RECT	3.515 51.53 3.565 51.66 ;
		RECT	4.51 51.53 4.56 51.66 ;
		RECT	5.035 51.53 5.085 51.66 ;
		RECT	6.22 51.53 6.27 51.66 ;
		RECT	7.5 51.53 7.55 51.66 ;
		RECT	9.72 51.53 9.77 51.66 ;
		RECT	11.025 51.53 11.075 51.66 ;
		RECT	13.8 52.21 13.85 52.34 ;
		RECT	3.02 52.66 3.15 52.71 ;
		RECT	1.57 52.685 1.62 52.815 ;
		RECT	4.87 52.685 4.92 52.815 ;
		RECT	6.375 52.685 6.425 52.815 ;
		RECT	7.015 52.685 7.065 52.815 ;
		RECT	10.27 52.685 10.32 52.815 ;
		RECT	12.79 52.685 12.84 52.815 ;
		RECT	14.33 52.685 14.38 52.815 ;
		RECT	3.02 52.79 3.15 52.84 ;
		RECT	4.035 53.18 4.085 53.31 ;
		RECT	12.655 53.18 12.705 53.31 ;
		RECT	13.9 53.18 13.95 53.31 ;
		RECT	3.02 53.65 3.15 53.7 ;
		RECT	1.57 53.675 1.62 53.805 ;
		RECT	4.87 53.675 4.92 53.805 ;
		RECT	6.375 53.675 6.425 53.805 ;
		RECT	7.015 53.675 7.065 53.805 ;
		RECT	10.27 53.675 10.32 53.805 ;
		RECT	12.79 53.675 12.84 53.805 ;
		RECT	14.33 53.675 14.38 53.805 ;
		RECT	3.02 53.78 3.15 53.83 ;
		RECT	0.62 54.165 0.67 54.295 ;
		RECT	3.65 54.165 3.7 54.295 ;
		RECT	7.19 54.165 7.24 54.295 ;
		RECT	14.14 54.165 14.19 54.295 ;
		RECT	6.85 54.45 6.9 54.5 ;
		RECT	1.045 54.63 1.175 54.68 ;
		RECT	1.34 54.63 1.47 54.68 ;
		RECT	4.47 54.63 4.6 54.68 ;
		RECT	1.86 54.655 1.91 54.785 ;
		RECT	2.01 54.655 2.06 54.785 ;
		RECT	2.32 54.655 2.37 54.785 ;
		RECT	3.25 54.655 3.3 54.785 ;
		RECT	3.515 54.655 3.565 54.785 ;
		RECT	5.035 54.655 5.085 54.785 ;
		RECT	6.22 54.655 6.27 54.785 ;
		RECT	7.5 54.655 7.55 54.785 ;
		RECT	9.72 54.655 9.77 54.785 ;
		RECT	11.025 54.655 11.075 54.785 ;
		RECT	1.045 54.76 1.175 54.81 ;
		RECT	1.34 54.76 1.47 54.81 ;
		RECT	4.47 54.76 4.6 54.81 ;
		RECT	0.9 55.125 14.055 55.305 ;
		RECT	3.02 55.615 3.15 55.665 ;
		RECT	1.57 55.64 1.62 55.77 ;
		RECT	4.87 55.64 4.92 55.77 ;
		RECT	6.375 55.64 6.425 55.77 ;
		RECT	7.015 55.64 7.065 55.77 ;
		RECT	10.27 55.64 10.32 55.77 ;
		RECT	12.79 55.64 12.84 55.77 ;
		RECT	14.33 55.64 14.38 55.77 ;
		RECT	3.02 55.745 3.15 55.795 ;
		RECT	4.035 56.135 4.085 56.265 ;
		RECT	12.655 56.135 12.705 56.265 ;
		RECT	13.9 56.135 13.95 56.265 ;
		RECT	3.02 56.6 3.15 56.65 ;
		RECT	1.57 56.625 1.62 56.755 ;
		RECT	4.87 56.625 4.92 56.755 ;
		RECT	6.375 56.625 6.425 56.755 ;
		RECT	7.015 56.625 7.065 56.755 ;
		RECT	10.27 56.625 10.32 56.755 ;
		RECT	12.79 56.625 12.84 56.755 ;
		RECT	14.33 56.625 14.38 56.755 ;
		RECT	3.02 56.73 3.15 56.78 ;
		RECT	6.85 56.91 6.9 56.96 ;
		RECT	4.035 57.115 4.085 57.245 ;
		RECT	12.655 57.115 12.705 57.245 ;
		RECT	3.02 57.585 3.15 57.635 ;
		RECT	1.57 57.61 1.62 57.74 ;
		RECT	4.87 57.61 4.92 57.74 ;
		RECT	6.375 57.61 6.425 57.74 ;
		RECT	10.27 57.61 10.32 57.74 ;
		RECT	12.79 57.61 12.84 57.74 ;
		RECT	14.33 57.61 14.38 57.74 ;
		RECT	3.02 57.715 3.15 57.765 ;
		RECT	3.8 58.075 3.93 58.125 ;
		RECT	5.635 58.075 5.765 58.125 ;
		RECT	8.31 58.075 8.44 58.125 ;
		RECT	8.73 58.075 8.86 58.125 ;
		RECT	0.9 58.1 0.95 58.23 ;
		RECT	2.485 58.1 2.535 58.23 ;
		RECT	2.615 58.1 2.665 58.23 ;
		RECT	6.065 58.1 6.115 58.23 ;
		RECT	6.725 58.1 6.775 58.23 ;
		RECT	11.555 58.1 12.57 58.23 ;
		RECT	14.005 58.1 14.055 58.23 ;
		RECT	3.8 58.205 3.93 58.255 ;
		RECT	5.635 58.205 5.765 58.255 ;
		RECT	8.31 58.205 8.44 58.255 ;
		RECT	8.73 58.205 8.86 58.255 ;
		RECT	1.045 58.57 1.175 58.62 ;
		RECT	1.34 58.57 1.47 58.62 ;
		RECT	4.47 58.57 4.6 58.62 ;
		RECT	9.275 58.57 9.405 58.62 ;
		RECT	1.86 58.595 1.91 58.725 ;
		RECT	2.01 58.595 2.06 58.725 ;
		RECT	2.32 58.595 2.37 58.725 ;
		RECT	3.25 58.595 3.3 58.725 ;
		RECT	3.515 58.595 3.565 58.725 ;
		RECT	6.22 58.595 6.27 58.725 ;
		RECT	7.5 58.595 7.55 58.725 ;
		RECT	9.72 58.595 9.77 58.725 ;
		RECT	11.025 58.595 11.075 58.725 ;
		RECT	1.045 58.7 1.175 58.75 ;
		RECT	1.34 58.7 1.47 58.75 ;
		RECT	4.47 58.7 4.6 58.75 ;
		RECT	9.275 58.7 9.405 58.75 ;
		RECT	3.8 59.06 3.93 59.11 ;
		RECT	5.635 59.06 5.765 59.11 ;
		RECT	8.31 59.06 8.44 59.11 ;
		RECT	8.73 59.06 8.86 59.11 ;
		RECT	0.9 59.085 0.95 59.215 ;
		RECT	2.485 59.085 2.535 59.215 ;
		RECT	2.615 59.085 2.665 59.215 ;
		RECT	6.065 59.085 6.115 59.215 ;
		RECT	6.725 59.085 6.775 59.215 ;
		RECT	11.555 59.085 11.865 59.215 ;
		RECT	12.52 59.085 12.57 59.215 ;
		RECT	14.005 59.085 14.055 59.215 ;
		RECT	3.8 59.19 3.93 59.24 ;
		RECT	5.635 59.19 5.765 59.24 ;
		RECT	8.31 59.19 8.44 59.24 ;
		RECT	8.73 59.19 8.86 59.24 ;
		RECT	3.02 59.55 3.15 59.6 ;
		RECT	1.57 59.575 1.62 59.705 ;
		RECT	4.87 59.575 4.92 59.705 ;
		RECT	6.375 59.575 6.425 59.705 ;
		RECT	10.27 59.575 10.32 59.705 ;
		RECT	12.79 59.575 12.84 59.705 ;
		RECT	14.33 59.575 14.38 59.705 ;
		RECT	3.02 59.68 3.15 59.73 ;
		RECT	0.9 60.045 14.055 60.225 ;
		RECT	3.02 60.535 3.15 60.585 ;
		RECT	1.57 60.56 1.62 60.69 ;
		RECT	4.87 60.56 4.92 60.69 ;
		RECT	6.375 60.56 6.425 60.69 ;
		RECT	10.27 60.56 10.32 60.69 ;
		RECT	12.79 60.56 12.84 60.69 ;
		RECT	14.33 60.56 14.38 60.69 ;
		RECT	3.02 60.665 3.15 60.715 ;
		RECT	12.655 61.045 12.705 61.175 ;
		RECT	4.035 61.055 4.085 61.185 ;
		RECT	3.02 61.52 3.15 61.57 ;
		RECT	1.57 61.545 1.62 61.675 ;
		RECT	4.87 61.545 4.92 61.675 ;
		RECT	6.375 61.545 6.425 61.675 ;
		RECT	10.27 61.545 10.32 61.675 ;
		RECT	12.79 61.545 12.84 61.675 ;
		RECT	14.33 61.545 14.38 61.675 ;
		RECT	3.02 61.65 3.15 61.7 ;
		RECT	0.9 62.01 14.055 62.19 ;
		RECT	14.29 62.32 14.42 62.37 ;
		RECT	1.045 62.505 1.175 62.555 ;
		RECT	1.34 62.505 1.47 62.555 ;
		RECT	4.47 62.505 4.6 62.555 ;
		RECT	9.275 62.505 9.405 62.555 ;
		RECT	1.86 62.53 1.91 62.66 ;
		RECT	2.01 62.53 2.06 62.66 ;
		RECT	2.32 62.53 2.37 62.66 ;
		RECT	3.25 62.53 3.3 62.66 ;
		RECT	3.515 62.53 3.565 62.66 ;
		RECT	6.22 62.53 6.27 62.66 ;
		RECT	7.5 62.53 7.55 62.66 ;
		RECT	9.72 62.53 9.77 62.66 ;
		RECT	11.025 62.53 11.075 62.66 ;
		RECT	1.045 62.635 1.175 62.685 ;
		RECT	1.34 62.635 1.47 62.685 ;
		RECT	4.47 62.635 4.6 62.685 ;
		RECT	9.275 62.635 9.405 62.685 ;
		RECT	0.9 62.815 0.95 62.865 ;
		RECT	2.51 62.815 2.64 62.865 ;
		RECT	0.9 62.995 14.055 63.175 ;
		RECT	2.18 63.515 2.23 63.645 ;
		RECT	8.56 63.515 8.61 63.645 ;
		RECT	10.27 63.515 10.32 63.645 ;
		RECT	4.035 64.005 4.085 64.135 ;
		RECT	3.02 64.47 3.15 64.52 ;
		RECT	1.57 64.495 1.62 64.625 ;
		RECT	4.87 64.495 4.92 64.625 ;
		RECT	6.375 64.495 6.425 64.625 ;
		RECT	11.69 64.495 11.74 64.625 ;
		RECT	12.79 64.495 12.84 64.625 ;
		RECT	12.79 64.495 12.84 64.625 ;
		RECT	14.33 64.495 14.38 64.625 ;
		RECT	3.02 64.6 3.15 64.65 ;
		RECT	4.035 64.955 4.085 65.085 ;
		RECT	12.655 64.955 12.705 65.085 ;
		RECT	3.02 65.455 3.15 65.505 ;
		RECT	1.57 65.48 1.62 65.61 ;
		RECT	4.87 65.48 4.92 65.61 ;
		RECT	6.375 65.48 6.425 65.61 ;
		RECT	11.69 65.48 11.74 65.61 ;
		RECT	12.79 65.48 12.84 65.61 ;
		RECT	12.79 65.48 12.84 65.61 ;
		RECT	14.33 65.48 14.38 65.61 ;
		RECT	3.02 65.585 3.15 65.635 ;
		RECT	0.9 65.915 14.055 66.095 ;
		RECT	1.045 66.455 1.175 66.505 ;
		RECT	1.34 66.455 1.47 66.505 ;
		RECT	4.47 66.455 4.6 66.505 ;
		RECT	9.275 66.455 9.405 66.505 ;
		RECT	1.86 66.48 1.91 66.61 ;
		RECT	2.01 66.48 2.06 66.61 ;
		RECT	3.25 66.48 3.3 66.61 ;
		RECT	3.515 66.48 3.565 66.61 ;
		RECT	6.22 66.48 6.27 66.61 ;
		RECT	7.5 66.48 7.55 66.61 ;
		RECT	9.72 66.48 9.77 66.61 ;
		RECT	11.025 66.48 11.075 66.61 ;
		RECT	1.045 66.585 1.175 66.635 ;
		RECT	1.34 66.585 1.47 66.635 ;
		RECT	4.47 66.585 4.6 66.635 ;
		RECT	9.275 66.585 9.405 66.635 ;
		RECT	12.655 66.755 12.705 66.805 ;
		RECT	1.045 66.93 1.175 66.98 ;
		RECT	1.34 66.93 1.47 66.98 ;
		RECT	4.47 66.93 4.6 66.98 ;
		RECT	9.275 66.93 9.405 66.98 ;
		RECT	1.86 66.955 1.91 67.085 ;
		RECT	2.01 66.955 2.06 67.085 ;
		RECT	3.25 66.955 3.3 67.085 ;
		RECT	3.515 66.955 3.565 67.085 ;
		RECT	6.22 66.955 6.27 67.085 ;
		RECT	7.5 66.955 7.55 67.085 ;
		RECT	9.72 66.955 9.77 67.085 ;
		RECT	11.025 66.955 11.075 67.085 ;
		RECT	13.675 66.955 13.725 67.085 ;
		RECT	1.045 67.06 1.175 67.11 ;
		RECT	1.34 67.06 1.47 67.11 ;
		RECT	4.47 67.06 4.6 67.11 ;
		RECT	9.275 67.06 9.405 67.11 ;
		RECT	3.02 67.425 3.15 67.475 ;
		RECT	1.57 67.45 1.62 67.58 ;
		RECT	4.87 67.45 4.92 67.58 ;
		RECT	6.375 67.45 6.425 67.58 ;
		RECT	8.975 67.45 9.025 67.58 ;
		RECT	11.69 67.45 11.74 67.58 ;
		RECT	12.79 67.45 12.84 67.58 ;
		RECT	14.33 67.45 14.38 67.58 ;
		RECT	3.02 67.555 3.15 67.605 ;
		RECT	12.655 67.735 12.705 67.785 ;
		RECT	0.9 67.915 14.055 68.095 ;
		RECT	1.57 68.435 1.62 68.565 ;
		RECT	4.87 68.435 4.92 68.565 ;
		RECT	6.375 68.435 6.425 68.565 ;
		RECT	8.975 68.435 9.025 68.565 ;
		RECT	11.69 68.435 11.74 68.565 ;
		RECT	12.79 68.435 12.84 68.565 ;
		RECT	14.33 68.435 14.38 68.565 ;
		RECT	3.02 68.475 3.15 68.525 ;
		RECT	1.045 68.72 1.175 68.77 ;
		RECT	1.34 68.72 1.47 68.77 ;
		RECT	4.47 68.72 4.6 68.77 ;
		RECT	9.275 68.72 9.405 68.77 ;
		RECT	1.86 68.745 1.91 68.875 ;
		RECT	2.01 68.745 2.06 68.875 ;
		RECT	3.25 68.745 3.3 68.875 ;
		RECT	3.515 68.745 3.565 68.875 ;
		RECT	6.22 68.745 6.27 68.875 ;
		RECT	7.5 68.745 7.55 68.875 ;
		RECT	9.72 68.745 9.77 68.875 ;
		RECT	11.025 68.745 11.075 68.875 ;
		RECT	1.045 68.85 1.175 68.9 ;
		RECT	1.34 68.85 1.47 68.9 ;
		RECT	4.47 68.85 4.6 68.9 ;
		RECT	9.275 68.85 9.405 68.9 ;
		RECT	13.8 69.225 13.85 69.355 ;
		RECT	2.18 69.455 2.23 69.585 ;
		RECT	8.56 69.455 8.61 69.585 ;
		RECT	10.27 69.455 10.32 69.585 ;
		RECT	0.62 69.685 0.67 69.815 ;
		RECT	3.65 69.685 3.7 69.815 ;
		RECT	7.19 69.685 7.24 69.815 ;
		RECT	14.14 69.685 14.19 69.815 ;
		RECT	1.085 69.915 1.135 70.045 ;
		RECT	1.38 69.915 1.43 70.045 ;
		RECT	1.86 69.915 1.91 70.045 ;
		RECT	2.01 69.915 2.06 70.045 ;
		RECT	3.25 69.915 3.3 70.045 ;
		RECT	3.515 69.915 3.565 70.045 ;
		RECT	4.51 69.915 4.56 70.045 ;
		RECT	6.22 69.915 6.27 70.045 ;
		RECT	7.5 69.915 7.55 70.045 ;
		RECT	9.315 69.915 9.365 70.045 ;
		RECT	9.72 69.915 9.77 70.045 ;
		RECT	11.025 69.915 11.075 70.045 ;
		RECT	0.435 29.565 0.485 29.695 ;
		RECT	0.435 30.545 0.485 30.675 ;
		RECT	0.435 32.515 0.485 32.645 ;
		RECT	0.435 33.5 0.485 33.63 ;
		RECT	0.435 36.455 0.485 36.585 ;
		RECT	0.435 37.435 0.485 37.565 ;
		RECT	0.435 38.42 0.485 38.55 ;
		RECT	0.435 40.39 0.485 40.52 ;
		RECT	0.17 41.17 0.22 41.22 ;
		RECT	0.435 41.37 0.485 41.5 ;
		RECT	0.435 42.355 0.485 42.485 ;
		RECT	0.18 43.135 0.23 43.185 ;
		RECT	0.435 44.33 0.485 44.46 ;
		RECT	0.435 45.31 0.485 45.44 ;
		RECT	0.435 48.26 0.485 48.39 ;
		RECT	0.435 49.735 0.485 49.865 ;
		RECT	0.435 52.685 0.485 52.815 ;
		RECT	0.435 53.675 0.485 53.805 ;
		RECT	0.18 54.45 0.23 54.5 ;
		RECT	0.435 55.64 0.485 55.77 ;
		RECT	0.435 56.625 0.485 56.755 ;
		RECT	0.17 56.91 0.22 56.96 ;
		RECT	0.435 57.61 0.485 57.74 ;
		RECT	0.435 59.575 0.485 59.705 ;
		RECT	0.435 60.56 0.485 60.69 ;
		RECT	0.435 61.545 0.485 61.675 ;
		RECT	0.17 62.815 0.22 62.865 ;
		RECT	0.435 63.8 0.485 63.85 ;
		RECT	0.435 64.29 0.485 64.34 ;
		RECT	0.435 64.495 0.485 64.625 ;
		RECT	0.435 65.48 0.485 65.61 ;
		RECT	0.435 67.45 0.485 67.58 ;
		RECT	0.435 68.435 0.485 68.565 ;
		RECT	3.06 69.915 3.11 70.045 ;
		RECT	4.87 69.915 4.92 70.045 ;
		RECT	6.375 69.915 6.425 70.045 ;
		RECT	8.975 69.915 9.025 70.045 ;
		RECT	12.79 69.915 12.84 70.045 ;
		RECT	1.57 28.015 1.62 28.145 ;
		RECT	3.06 28.015 3.11 28.145 ;
		RECT	4.87 28.015 4.92 28.145 ;
		RECT	12.79 28.015 12.84 28.145 ;
		RECT	1.57 29.18 1.62 29.31 ;
		RECT	3.02 29.155 3.15 29.335 ;
		RECT	4.87 29.18 4.92 29.31 ;
		RECT	8.955 29.18 9.005 29.31 ;
		RECT	12.79 29.18 12.84 29.31 ;
		RECT	14.29 29.155 14.42 29.335 ;
		RECT	1.045 29.54 1.175 29.72 ;
		RECT	1.34 29.54 1.47 29.72 ;
		RECT	1.86 29.565 1.91 29.695 ;
		RECT	2.01 29.565 2.06 29.695 ;
		RECT	3.25 29.565 3.3 29.695 ;
		RECT	3.515 29.565 3.565 29.695 ;
		RECT	4.47 29.54 4.6 29.72 ;
		RECT	5.035 29.565 5.085 29.695 ;
		RECT	6.22 29.565 6.27 29.695 ;
		RECT	7.5 29.565 7.55 29.695 ;
		RECT	9.275 29.54 9.405 29.72 ;
		RECT	9.72 29.565 9.77 29.695 ;
		RECT	11.025 29.565 11.075 29.695 ;
		RECT	1.045 30.52 1.175 30.7 ;
		RECT	1.34 30.52 1.47 30.7 ;
		RECT	1.86 30.545 1.91 30.675 ;
		RECT	2.01 30.545 2.06 30.675 ;
		RECT	3.25 30.545 3.3 30.675 ;
		RECT	3.515 30.545 3.565 30.675 ;
		RECT	4.47 30.52 4.6 30.7 ;
		RECT	5.035 30.545 5.085 30.675 ;
		RECT	6.22 30.545 6.27 30.675 ;
		RECT	7.5 30.545 7.55 30.675 ;
		RECT	9.275 30.52 9.405 30.7 ;
		RECT	9.72 30.545 9.77 30.675 ;
		RECT	11.025 30.545 11.075 30.675 ;
		RECT	1.57 31.045 1.62 31.175 ;
		RECT	3.02 31.02 3.15 31.2 ;
		RECT	4.87 31.045 4.92 31.175 ;
		RECT	5.9 31.045 5.95 31.175 ;
		RECT	8.955 31.045 9.005 31.175 ;
		RECT	1.57 31.515 1.62 31.645 ;
		RECT	3.02 31.49 3.15 31.67 ;
		RECT	4.87 31.515 4.92 31.645 ;
		RECT	5.9 31.515 5.95 31.645 ;
		RECT	8.955 31.515 9.005 31.645 ;
		RECT	12.79 31.515 12.84 31.645 ;
		RECT	1.045 32.49 1.175 32.67 ;
		RECT	1.34 32.49 1.47 32.67 ;
		RECT	1.86 32.515 1.91 32.645 ;
		RECT	2.01 32.515 2.06 32.645 ;
		RECT	3.25 32.515 3.3 32.645 ;
		RECT	3.515 32.515 3.565 32.645 ;
		RECT	4.47 32.49 4.6 32.67 ;
		RECT	5.035 32.515 5.085 32.645 ;
		RECT	6.22 32.515 6.27 32.645 ;
		RECT	7.5 32.515 7.55 32.645 ;
		RECT	9.275 32.49 9.405 32.67 ;
		RECT	9.72 32.515 9.77 32.645 ;
		RECT	11.025 32.515 11.075 32.645 ;
		RECT	1.045 33.475 1.175 33.655 ;
		RECT	1.34 33.475 1.47 33.655 ;
		RECT	1.86 33.5 1.91 33.63 ;
		RECT	2.01 33.5 2.06 33.63 ;
		RECT	3.25 33.5 3.3 33.63 ;
		RECT	3.515 33.5 3.565 33.63 ;
		RECT	4.47 33.475 4.6 33.655 ;
		RECT	5.035 33.5 5.085 33.63 ;
		RECT	6.22 33.5 6.27 33.63 ;
		RECT	7.5 33.5 7.55 33.63 ;
		RECT	9.72 33.5 9.77 33.63 ;
		RECT	11.025 33.5 11.075 33.63 ;
		RECT	1.57 35.47 1.62 35.6 ;
		RECT	3.02 35.445 3.15 35.625 ;
		RECT	4.87 35.47 4.92 35.6 ;
		RECT	5.9 35.47 5.95 35.6 ;
		RECT	12.79 35.47 12.84 35.6 ;
		RECT	14.29 35.445 14.42 35.625 ;
		RECT	1.045 36.43 1.175 36.61 ;
		RECT	1.34 36.43 1.47 36.61 ;
		RECT	1.86 36.455 1.91 36.585 ;
		RECT	2.01 36.455 2.06 36.585 ;
		RECT	2.32 36.455 2.37 36.585 ;
		RECT	3.25 36.455 3.3 36.585 ;
		RECT	3.515 36.455 3.565 36.585 ;
		RECT	4.47 36.43 4.6 36.61 ;
		RECT	5.035 36.455 5.085 36.585 ;
		RECT	6.22 36.455 6.27 36.585 ;
		RECT	7.5 36.455 7.55 36.585 ;
		RECT	9.72 36.455 9.77 36.585 ;
		RECT	11.025 36.455 11.075 36.585 ;
		RECT	1.045 37.41 1.175 37.59 ;
		RECT	1.34 37.41 1.47 37.59 ;
		RECT	1.86 37.435 1.91 37.565 ;
		RECT	2.01 37.435 2.06 37.565 ;
		RECT	2.32 37.435 2.37 37.565 ;
		RECT	3.25 37.435 3.3 37.565 ;
		RECT	3.515 37.435 3.565 37.565 ;
		RECT	4.47 37.41 4.6 37.59 ;
		RECT	5.035 37.435 5.085 37.565 ;
		RECT	6.22 37.435 6.27 37.565 ;
		RECT	7.5 37.435 7.55 37.565 ;
		RECT	9.72 37.435 9.77 37.565 ;
		RECT	11.025 37.435 11.075 37.565 ;
		RECT	1.045 38.395 1.175 38.575 ;
		RECT	1.34 38.395 1.47 38.575 ;
		RECT	1.86 38.42 1.91 38.55 ;
		RECT	2.01 38.42 2.06 38.55 ;
		RECT	2.32 38.42 2.37 38.55 ;
		RECT	3.25 38.42 3.3 38.55 ;
		RECT	3.515 38.42 3.565 38.55 ;
		RECT	4.47 38.395 4.6 38.575 ;
		RECT	5.035 38.42 5.085 38.55 ;
		RECT	6.22 38.42 6.27 38.55 ;
		RECT	7.5 38.42 7.55 38.55 ;
		RECT	9.72 38.42 9.77 38.55 ;
		RECT	11.025 38.42 11.075 38.55 ;
		RECT	1.57 39.405 1.62 39.535 ;
		RECT	3.02 39.38 3.15 39.56 ;
		RECT	4.87 39.405 4.92 39.535 ;
		RECT	5.9 39.405 5.95 39.535 ;
		RECT	9.43 39.405 9.48 39.535 ;
		RECT	10.27 39.405 10.32 39.535 ;
		RECT	12.79 39.405 12.84 39.535 ;
		RECT	14.29 39.38 14.42 39.56 ;
		RECT	1.045 40.365 1.175 40.545 ;
		RECT	1.34 40.365 1.47 40.545 ;
		RECT	1.86 40.39 1.91 40.52 ;
		RECT	2.01 40.39 2.06 40.52 ;
		RECT	2.32 40.39 2.37 40.52 ;
		RECT	3.25 40.39 3.3 40.52 ;
		RECT	3.515 40.39 3.565 40.52 ;
		RECT	4.47 40.365 4.6 40.545 ;
		RECT	5.035 40.39 5.085 40.52 ;
		RECT	6.22 40.39 6.27 40.52 ;
		RECT	7.5 40.39 7.55 40.52 ;
		RECT	9.72 40.39 9.77 40.52 ;
		RECT	11.025 40.39 11.075 40.52 ;
		RECT	1.045 41.345 1.175 41.525 ;
		RECT	1.34 41.345 1.47 41.525 ;
		RECT	1.86 41.37 1.91 41.5 ;
		RECT	2.01 41.37 2.06 41.5 ;
		RECT	2.32 41.37 2.37 41.5 ;
		RECT	3.25 41.37 3.3 41.5 ;
		RECT	3.515 41.37 3.565 41.5 ;
		RECT	4.47 41.345 4.6 41.525 ;
		RECT	5.035 41.37 5.085 41.5 ;
		RECT	6.22 41.37 6.27 41.5 ;
		RECT	7.5 41.37 7.55 41.5 ;
		RECT	9.72 41.37 9.77 41.5 ;
		RECT	11.025 41.37 11.075 41.5 ;
		RECT	1.045 42.33 1.175 42.51 ;
		RECT	1.34 42.33 1.47 42.51 ;
		RECT	1.86 42.355 1.91 42.485 ;
		RECT	2.01 42.355 2.06 42.485 ;
		RECT	2.32 42.355 2.37 42.485 ;
		RECT	3.25 42.355 3.3 42.485 ;
		RECT	3.515 42.355 3.565 42.485 ;
		RECT	4.47 42.33 4.6 42.51 ;
		RECT	5.035 42.355 5.085 42.485 ;
		RECT	6.22 42.355 6.27 42.485 ;
		RECT	7.5 42.355 7.55 42.485 ;
		RECT	9.72 42.355 9.77 42.485 ;
		RECT	11.025 42.355 11.075 42.485 ;
		RECT	1.57 43.34 1.62 43.47 ;
		RECT	3.02 43.315 3.15 43.495 ;
		RECT	4.87 43.34 4.92 43.47 ;
		RECT	5.9 43.34 5.95 43.47 ;
		RECT	6.375 43.34 6.425 43.47 ;
		RECT	7.015 43.34 7.065 43.47 ;
		RECT	10.27 43.34 10.32 43.47 ;
		RECT	12.79 43.34 12.84 43.47 ;
		RECT	14.29 43.315 14.42 43.495 ;
		RECT	1.045 44.305 1.175 44.485 ;
		RECT	1.34 44.305 1.47 44.485 ;
		RECT	1.86 44.33 1.91 44.46 ;
		RECT	2.01 44.33 2.06 44.46 ;
		RECT	2.32 44.33 2.37 44.46 ;
		RECT	3.25 44.33 3.3 44.46 ;
		RECT	3.515 44.33 3.565 44.46 ;
		RECT	4.47 44.305 4.6 44.485 ;
		RECT	5.035 44.33 5.085 44.46 ;
		RECT	6.22 44.33 6.27 44.46 ;
		RECT	7.5 44.33 7.55 44.46 ;
		RECT	9.72 44.33 9.77 44.46 ;
		RECT	11.025 44.33 11.075 44.46 ;
		RECT	1.045 45.285 1.175 45.465 ;
		RECT	1.34 45.285 1.47 45.465 ;
		RECT	1.86 45.31 1.91 45.44 ;
		RECT	2.01 45.31 2.06 45.44 ;
		RECT	2.32 45.31 2.37 45.44 ;
		RECT	3.25 45.31 3.3 45.44 ;
		RECT	3.515 45.31 3.565 45.44 ;
		RECT	4.47 45.285 4.6 45.465 ;
		RECT	5.035 45.31 5.085 45.44 ;
		RECT	6.22 45.31 6.27 45.44 ;
		RECT	7.5 45.31 7.55 45.44 ;
		RECT	9.72 45.31 9.77 45.44 ;
		RECT	11.025 45.31 11.075 45.44 ;
		RECT	1.57 46.465 1.62 46.595 ;
		RECT	3.06 46.465 3.11 46.595 ;
		RECT	4.87 46.465 4.92 46.595 ;
		RECT	5.9 46.465 5.95 46.595 ;
		RECT	6.375 46.465 6.425 46.595 ;
		RECT	7.015 46.465 7.065 46.595 ;
		RECT	9.11 46.465 9.16 46.595 ;
		RECT	10.27 46.465 10.32 46.595 ;
		RECT	1.57 47.275 1.62 47.405 ;
		RECT	3.02 47.25 3.15 47.43 ;
		RECT	4.87 47.275 4.92 47.405 ;
		RECT	5.9 47.275 5.95 47.405 ;
		RECT	6.375 47.275 6.425 47.405 ;
		RECT	7.015 47.275 7.065 47.405 ;
		RECT	9.11 47.275 9.16 47.405 ;
		RECT	10.27 47.275 10.32 47.405 ;
		RECT	12.79 47.275 12.84 47.405 ;
		RECT	1.045 48.235 1.175 48.415 ;
		RECT	1.34 48.235 1.47 48.415 ;
		RECT	1.86 48.26 1.91 48.39 ;
		RECT	2.01 48.26 2.06 48.39 ;
		RECT	2.32 48.26 2.37 48.39 ;
		RECT	3.25 48.26 3.3 48.39 ;
		RECT	3.515 48.26 3.565 48.39 ;
		RECT	4.47 48.235 4.6 48.415 ;
		RECT	5.035 48.26 5.085 48.39 ;
		RECT	6.22 48.26 6.27 48.39 ;
		RECT	7.5 48.26 7.55 48.39 ;
		RECT	9.72 48.26 9.77 48.39 ;
		RECT	11.025 48.26 11.075 48.39 ;
		RECT	1.045 49.71 1.175 49.89 ;
		RECT	1.34 49.71 1.47 49.89 ;
		RECT	1.86 49.735 1.91 49.865 ;
		RECT	2.01 49.735 2.06 49.865 ;
		RECT	2.32 49.735 2.37 49.865 ;
		RECT	3.25 49.735 3.3 49.865 ;
		RECT	3.515 49.735 3.565 49.865 ;
		RECT	4.47 49.71 4.6 49.89 ;
		RECT	5.035 49.735 5.085 49.865 ;
		RECT	6.22 49.735 6.27 49.865 ;
		RECT	7.5 49.735 7.55 49.865 ;
		RECT	9.72 49.735 9.77 49.865 ;
		RECT	11.025 49.735 11.075 49.865 ;
		RECT	1.57 50.72 1.62 50.85 ;
		RECT	3.02 50.695 3.15 50.875 ;
		RECT	4.87 50.72 4.92 50.85 ;
		RECT	6.375 50.72 6.425 50.85 ;
		RECT	7.015 50.72 7.065 50.85 ;
		RECT	9.11 50.72 9.16 50.85 ;
		RECT	10.27 50.72 10.32 50.85 ;
		RECT	12.79 50.72 12.84 50.85 ;
		RECT	1.57 51.53 1.62 51.66 ;
		RECT	3.06 51.53 3.11 51.66 ;
		RECT	4.87 51.53 4.92 51.66 ;
		RECT	6.375 51.53 6.425 51.66 ;
		RECT	7.015 51.53 7.065 51.66 ;
		RECT	9.11 51.53 9.16 51.66 ;
		RECT	10.27 51.53 10.32 51.66 ;
		RECT	1.045 52.66 1.175 52.84 ;
		RECT	1.34 52.66 1.47 52.84 ;
		RECT	1.86 52.685 1.91 52.815 ;
		RECT	2.01 52.685 2.06 52.815 ;
		RECT	2.32 52.685 2.37 52.815 ;
		RECT	3.25 52.685 3.3 52.815 ;
		RECT	3.515 52.685 3.565 52.815 ;
		RECT	4.47 52.66 4.6 52.84 ;
		RECT	5.035 52.685 5.085 52.815 ;
		RECT	6.22 52.685 6.27 52.815 ;
		RECT	7.5 52.685 7.55 52.815 ;
		RECT	9.72 52.685 9.77 52.815 ;
		RECT	11.025 52.685 11.075 52.815 ;
		RECT	1.045 53.65 1.175 53.83 ;
		RECT	1.34 53.65 1.47 53.83 ;
		RECT	1.86 53.675 1.91 53.805 ;
		RECT	2.01 53.675 2.06 53.805 ;
		RECT	2.32 53.675 2.37 53.805 ;
		RECT	3.25 53.675 3.3 53.805 ;
		RECT	3.515 53.675 3.565 53.805 ;
		RECT	4.47 53.65 4.6 53.83 ;
		RECT	5.035 53.675 5.085 53.805 ;
		RECT	6.22 53.675 6.27 53.805 ;
		RECT	7.5 53.675 7.55 53.805 ;
		RECT	9.72 53.675 9.77 53.805 ;
		RECT	11.025 53.675 11.075 53.805 ;
		RECT	1.57 54.655 1.62 54.785 ;
		RECT	3.02 54.63 3.15 54.81 ;
		RECT	4.87 54.655 4.92 54.785 ;
		RECT	6.375 54.655 6.425 54.785 ;
		RECT	7.015 54.655 7.065 54.785 ;
		RECT	10.27 54.655 10.32 54.785 ;
		RECT	12.79 54.655 12.84 54.785 ;
		RECT	14.29 54.63 14.42 54.81 ;
		RECT	1.045 55.615 1.175 55.795 ;
		RECT	1.34 55.615 1.47 55.795 ;
		RECT	1.86 55.64 1.91 55.77 ;
		RECT	2.01 55.64 2.06 55.77 ;
		RECT	2.32 55.64 2.37 55.77 ;
		RECT	3.25 55.64 3.3 55.77 ;
		RECT	3.515 55.64 3.565 55.77 ;
		RECT	4.47 55.615 4.6 55.795 ;
		RECT	5.035 55.64 5.085 55.77 ;
		RECT	6.22 55.64 6.27 55.77 ;
		RECT	7.5 55.64 7.55 55.77 ;
		RECT	9.275 55.615 9.405 55.795 ;
		RECT	9.72 55.64 9.77 55.77 ;
		RECT	11.025 55.64 11.075 55.77 ;
		RECT	1.045 56.6 1.175 56.78 ;
		RECT	1.34 56.6 1.47 56.78 ;
		RECT	1.86 56.625 1.91 56.755 ;
		RECT	2.01 56.625 2.06 56.755 ;
		RECT	2.32 56.625 2.37 56.755 ;
		RECT	3.25 56.625 3.3 56.755 ;
		RECT	3.515 56.625 3.565 56.755 ;
		RECT	4.47 56.6 4.6 56.78 ;
		RECT	5.035 56.625 5.085 56.755 ;
		RECT	6.22 56.625 6.27 56.755 ;
		RECT	7.5 56.625 7.55 56.755 ;
		RECT	9.275 56.6 9.405 56.78 ;
		RECT	9.72 56.625 9.77 56.755 ;
		RECT	11.025 56.625 11.075 56.755 ;
		RECT	1.045 57.585 1.175 57.765 ;
		RECT	1.34 57.585 1.47 57.765 ;
		RECT	1.86 57.61 1.91 57.74 ;
		RECT	2.01 57.61 2.06 57.74 ;
		RECT	2.32 57.61 2.37 57.74 ;
		RECT	3.25 57.61 3.3 57.74 ;
		RECT	3.515 57.61 3.565 57.74 ;
		RECT	4.47 57.585 4.6 57.765 ;
		RECT	6.22 57.61 6.27 57.74 ;
		RECT	7.5 57.61 7.55 57.74 ;
		RECT	9.275 57.585 9.405 57.765 ;
		RECT	9.72 57.61 9.77 57.74 ;
		RECT	11.025 57.61 11.075 57.74 ;
		RECT	1.57 58.595 1.62 58.725 ;
		RECT	3.02 58.57 3.15 58.75 ;
		RECT	4.87 58.595 4.92 58.725 ;
		RECT	6.375 58.595 6.425 58.725 ;
		RECT	10 58.595 10.05 58.725 ;
		RECT	10.27 58.595 10.32 58.725 ;
		RECT	12.79 58.595 12.84 58.725 ;
		RECT	14.29 58.57 14.42 58.75 ;
		RECT	1.045 59.55 1.175 59.73 ;
		RECT	1.34 59.55 1.47 59.73 ;
		RECT	1.86 59.575 1.91 59.705 ;
		RECT	2.01 59.575 2.06 59.705 ;
		RECT	2.32 59.575 2.37 59.705 ;
		RECT	3.25 59.575 3.3 59.705 ;
		RECT	3.515 59.575 3.565 59.705 ;
		RECT	4.47 59.55 4.6 59.73 ;
		RECT	6.22 59.575 6.27 59.705 ;
		RECT	7.5 59.575 7.55 59.705 ;
		RECT	9.275 59.55 9.405 59.73 ;
		RECT	9.72 59.575 9.77 59.705 ;
		RECT	11.025 59.575 11.075 59.705 ;
		RECT	1.045 60.535 1.175 60.715 ;
		RECT	1.34 60.535 1.47 60.715 ;
		RECT	1.86 60.56 1.91 60.69 ;
		RECT	2.01 60.56 2.06 60.69 ;
		RECT	2.32 60.56 2.37 60.69 ;
		RECT	3.25 60.56 3.3 60.69 ;
		RECT	3.515 60.56 3.565 60.69 ;
		RECT	4.47 60.535 4.6 60.715 ;
		RECT	6.22 60.56 6.27 60.69 ;
		RECT	7.5 60.56 7.55 60.69 ;
		RECT	9.275 60.535 9.405 60.715 ;
		RECT	9.72 60.56 9.77 60.69 ;
		RECT	11.025 60.56 11.075 60.69 ;
		RECT	1.045 61.52 1.175 61.7 ;
		RECT	1.34 61.52 1.47 61.7 ;
		RECT	1.86 61.545 1.91 61.675 ;
		RECT	2.01 61.545 2.06 61.675 ;
		RECT	2.32 61.545 2.37 61.675 ;
		RECT	3.25 61.545 3.3 61.675 ;
		RECT	3.515 61.545 3.565 61.675 ;
		RECT	4.47 61.52 4.6 61.7 ;
		RECT	6.22 61.545 6.27 61.675 ;
		RECT	7.5 61.545 7.55 61.675 ;
		RECT	9.275 61.52 9.405 61.7 ;
		RECT	9.72 61.545 9.77 61.675 ;
		RECT	11.025 61.545 11.075 61.675 ;
		RECT	1.57 62.53 1.62 62.66 ;
		RECT	3.02 62.505 3.15 62.685 ;
		RECT	4.87 62.53 4.92 62.66 ;
		RECT	6.375 62.53 6.425 62.66 ;
		RECT	12.79 62.53 12.84 62.66 ;
		RECT	14.29 62.505 14.42 62.685 ;
		RECT	1.045 64.47 1.175 64.65 ;
		RECT	1.34 64.47 1.47 64.65 ;
		RECT	1.86 64.495 1.91 64.625 ;
		RECT	2.01 64.495 2.06 64.625 ;
		RECT	2.32 64.495 2.37 64.625 ;
		RECT	3.25 64.495 3.3 64.625 ;
		RECT	3.515 64.495 3.565 64.625 ;
		RECT	4.47 64.47 4.6 64.65 ;
		RECT	6.22 64.495 6.27 64.625 ;
		RECT	7.5 64.495 7.55 64.625 ;
		RECT	9.275 64.47 9.405 64.65 ;
		RECT	9.72 64.495 9.77 64.625 ;
		RECT	11.025 64.495 11.075 64.625 ;
		RECT	1.045 65.455 1.175 65.635 ;
		RECT	1.34 65.455 1.47 65.635 ;
		RECT	1.86 65.48 1.91 65.61 ;
		RECT	2.01 65.48 2.06 65.61 ;
		RECT	2.32 65.48 2.37 65.61 ;
		RECT	3.25 65.48 3.3 65.61 ;
		RECT	3.515 65.48 3.565 65.61 ;
		RECT	4.47 65.455 4.6 65.635 ;
		RECT	6.22 65.48 6.27 65.61 ;
		RECT	7.5 65.48 7.55 65.61 ;
		RECT	9.275 65.455 9.405 65.635 ;
		RECT	9.72 65.48 9.77 65.61 ;
		RECT	11.025 65.48 11.075 65.61 ;
		RECT	1.57 66.48 1.62 66.61 ;
		RECT	3.02 66.455 3.15 66.635 ;
		RECT	4.87 66.48 4.92 66.61 ;
		RECT	6.375 66.48 6.425 66.61 ;
		RECT	11.69 66.48 11.74 66.61 ;
		RECT	12.79 66.48 12.84 66.61 ;
		RECT	1.57 66.955 1.62 67.085 ;
		RECT	3.02 66.93 3.15 67.11 ;
		RECT	4.87 66.955 4.92 67.085 ;
		RECT	6.375 66.955 6.425 67.085 ;
		RECT	1.045 67.425 1.175 67.605 ;
		RECT	1.34 67.425 1.47 67.605 ;
		RECT	1.86 67.45 1.91 67.58 ;
		RECT	2.01 67.45 2.06 67.58 ;
		RECT	3.25 67.45 3.3 67.58 ;
		RECT	3.515 67.45 3.565 67.58 ;
		RECT	4.47 67.425 4.6 67.605 ;
		RECT	6.22 67.45 6.27 67.58 ;
		RECT	7.5 67.45 7.55 67.58 ;
		RECT	9.275 67.425 9.405 67.605 ;
		RECT	9.72 67.45 9.77 67.58 ;
		RECT	11.025 67.45 11.075 67.58 ;
		RECT	1.86 68.435 1.91 68.565 ;
		RECT	2.01 68.435 2.06 68.565 ;
		RECT	3.25 68.435 3.3 68.565 ;
		RECT	3.515 68.435 3.565 68.565 ;
		RECT	6.22 68.435 6.27 68.565 ;
		RECT	7.5 68.435 7.55 68.565 ;
		RECT	9.72 68.435 9.77 68.565 ;
		RECT	11.025 68.435 11.075 68.565 ;
		RECT	1.57 68.745 1.62 68.875 ;
		RECT	3.02 68.72 3.15 68.9 ;
		RECT	4.87 68.745 4.92 68.875 ;
		RECT	6.375 68.745 6.425 68.875 ;
		RECT	8.975 68.745 9.025 68.875 ;
		RECT	12.79 68.745 12.84 68.875 ;
		RECT	14.29 68.72 14.42 68.9 ;
		RECT	0.9 28.245 0.95 28.375 ;
		RECT	2.485 28.245 2.665 28.375 ;
		RECT	3.84 28.245 3.89 28.375 ;
		RECT	5.675 28.245 5.725 28.375 ;
		RECT	6.065 28.245 6.115 28.375 ;
		RECT	6.725 28.245 6.775 28.375 ;
		RECT	8.35 28.245 8.4 28.375 ;
		RECT	8.77 28.245 8.82 28.375 ;
		RECT	11.555 28.245 11.605 28.375 ;
		RECT	11.815 28.245 11.865 28.375 ;
		RECT	12.52 28.245 12.57 28.375 ;
		RECT	14.005 28.245 14.055 28.375 ;
		RECT	0.62 30.055 0.67 30.185 ;
		RECT	3.65 30.055 3.7 30.185 ;
		RECT	7.18 30.055 7.23 30.185 ;
		RECT	14.14 30.055 14.19 30.185 ;
		RECT	0.62 32.06 0.67 32.19 ;
		RECT	3.65 32.06 3.7 32.19 ;
		RECT	7.18 32.06 7.23 32.19 ;
		RECT	14.14 32.06 14.19 32.19 ;
		RECT	0.62 34.975 0.67 35.105 ;
		RECT	3.65 34.975 3.7 35.105 ;
		RECT	7.18 34.975 7.23 35.105 ;
		RECT	14.14 34.975 14.19 35.105 ;
		RECT	0.62 35.96 0.67 36.09 ;
		RECT	3.65 35.96 3.7 36.09 ;
		RECT	7.18 35.96 7.23 36.09 ;
		RECT	14.14 35.96 14.19 36.09 ;
		RECT	0.62 37.93 0.67 38.06 ;
		RECT	3.65 37.93 3.7 38.06 ;
		RECT	7.18 37.93 7.23 38.06 ;
		RECT	14.14 37.93 14.19 38.06 ;
		RECT	0.62 38.91 0.67 39.04 ;
		RECT	3.65 38.91 3.7 39.04 ;
		RECT	7.18 38.91 7.23 39.04 ;
		RECT	14.14 38.91 14.19 39.04 ;
		RECT	0.62 39.895 0.67 40.025 ;
		RECT	3.65 39.895 3.7 40.025 ;
		RECT	7.18 39.895 7.23 40.025 ;
		RECT	14.14 39.895 14.19 40.025 ;
		RECT	0.62 42.85 0.67 42.98 ;
		RECT	3.65 42.85 3.7 42.98 ;
		RECT	7.18 42.85 7.23 42.98 ;
		RECT	14.14 42.85 14.19 42.98 ;
		RECT	0.9 43.835 0.95 43.965 ;
		RECT	2.485 43.835 2.665 43.965 ;
		RECT	3.8 43.81 3.93 43.99 ;
		RECT	5.635 43.81 5.765 43.99 ;
		RECT	6.065 43.835 6.115 43.965 ;
		RECT	6.675 43.835 6.725 43.965 ;
		RECT	8.31 43.81 8.44 43.99 ;
		RECT	8.73 43.81 8.86 43.99 ;
		RECT	11.555 43.835 11.605 43.965 ;
		RECT	11.815 43.835 11.865 43.965 ;
		RECT	12.52 43.835 12.57 43.965 ;
		RECT	14.005 43.835 14.055 43.965 ;
		RECT	0.62 46.785 0.67 46.915 ;
		RECT	3.65 46.785 3.7 46.915 ;
		RECT	7.18 46.785 7.23 46.915 ;
		RECT	14.14 46.785 14.19 46.915 ;
		RECT	0.62 47.77 0.67 47.9 ;
		RECT	3.65 47.77 3.7 47.9 ;
		RECT	7.18 47.77 7.23 47.9 ;
		RECT	14.14 47.77 14.19 47.9 ;
		RECT	8.31 49.04 8.44 49.09 ;
		RECT	8.73 49.04 8.86 49.09 ;
		RECT	10.12 49.04 10.17 49.09 ;
		RECT	11.555 49.04 11.605 49.09 ;
		RECT	11.815 49.04 11.865 49.09 ;
		RECT	12.52 49.04 12.57 49.09 ;
		RECT	0.62 50.23 0.67 50.36 ;
		RECT	3.65 50.23 3.7 50.36 ;
		RECT	7.18 50.23 7.23 50.36 ;
		RECT	12.655 50.23 12.705 50.36 ;
		RECT	14.14 50.23 14.19 50.36 ;
		RECT	0.62 51.21 0.67 51.34 ;
		RECT	3.65 51.21 3.7 51.34 ;
		RECT	7.18 51.21 7.23 51.34 ;
		RECT	14.14 51.21 14.19 51.34 ;
		RECT	0.9 54.165 0.95 54.295 ;
		RECT	2.51 54.14 2.64 54.32 ;
		RECT	3.8 54.14 3.93 54.32 ;
		RECT	5.635 54.14 5.765 54.32 ;
		RECT	6.065 54.165 6.115 54.295 ;
		RECT	6.675 54.165 6.725 54.295 ;
		RECT	8.31 54.14 8.44 54.32 ;
		RECT	8.73 54.14 8.86 54.32 ;
		RECT	11.555 54.165 11.605 54.295 ;
		RECT	11.815 54.165 11.865 54.295 ;
		RECT	12.52 54.165 12.57 54.295 ;
		RECT	14.005 54.165 14.055 54.295 ;
		RECT	0.62 55.15 0.67 55.28 ;
		RECT	3.65 55.15 3.7 55.28 ;
		RECT	7.18 55.15 7.23 55.28 ;
		RECT	14.14 55.15 14.19 55.28 ;
		RECT	0.62 58.1 0.67 58.23 ;
		RECT	3.65 58.1 3.7 58.23 ;
		RECT	7.18 58.1 7.23 58.23 ;
		RECT	14.14 58.1 14.19 58.23 ;
		RECT	0.62 59.085 0.67 59.215 ;
		RECT	3.65 59.085 3.7 59.215 ;
		RECT	7.18 59.085 7.23 59.215 ;
		RECT	14.14 59.085 14.19 59.215 ;
		RECT	0.62 60.07 0.67 60.2 ;
		RECT	3.65 60.07 3.7 60.2 ;
		RECT	7.18 60.07 7.23 60.2 ;
		RECT	14.14 60.07 14.19 60.2 ;
		RECT	0.62 62.035 0.67 62.165 ;
		RECT	3.65 62.035 3.7 62.165 ;
		RECT	7.18 62.035 7.23 62.165 ;
		RECT	14.14 62.035 14.19 62.165 ;
		RECT	0.62 62.815 0.67 62.865 ;
		RECT	0.62 63.02 0.67 63.15 ;
		RECT	3.65 63.02 3.7 63.15 ;
		RECT	7.18 63.02 7.23 63.15 ;
		RECT	14.14 63.02 14.19 63.15 ;
		RECT	0.62 65.94 0.67 66.07 ;
		RECT	3.65 65.94 3.7 66.07 ;
		RECT	7.18 65.94 7.23 66.07 ;
		RECT	14.14 65.94 14.19 66.07 ;
		RECT	0.62 67.94 0.67 68.07 ;
		RECT	3.65 67.94 3.7 68.07 ;
		RECT	7.18 67.94 7.23 68.07 ;
		RECT	14.14 67.94 14.19 68.07 ;
		RECT	0.9 69.685 0.95 69.815 ;
		RECT	2.485 69.685 2.665 69.815 ;
		RECT	3.84 69.685 3.89 69.815 ;
		RECT	5.675 69.685 5.725 69.815 ;
		RECT	6.065 69.685 6.115 69.815 ;
		RECT	6.725 69.685 6.775 69.815 ;
		RECT	8.35 69.685 8.4 69.815 ;
		RECT	8.77 69.685 8.82 69.815 ;
		RECT	11.555 69.685 11.605 69.815 ;
		RECT	11.815 69.685 11.865 69.815 ;
		RECT	12.52 69.685 12.57 69.815 ;
		RECT	14.005 69.685 14.055 69.815 ;
		RECT	1.57 28.475 1.62 28.605 ;
		RECT	3.06 28.475 3.11 28.605 ;
		RECT	4.87 28.475 4.92 28.605 ;
		RECT	12.79 28.475 12.84 28.605 ;
		RECT	14.33 28.475 14.38 28.605 ;
		RECT	2.18 29.565 2.23 29.695 ;
		RECT	8.56 29.565 8.61 29.695 ;
		RECT	10.27 29.565 10.32 29.695 ;
		RECT	2.18 30.545 2.23 30.675 ;
		RECT	8.56 30.545 8.61 30.675 ;
		RECT	10.27 30.545 10.32 30.675 ;
		RECT	2.18 32.515 2.23 32.645 ;
		RECT	8.56 32.515 8.61 32.645 ;
		RECT	10.27 32.515 10.32 32.645 ;
		RECT	2.18 33.5 2.23 33.63 ;
		RECT	8.56 33.5 8.61 33.63 ;
		RECT	10.27 33.5 10.32 33.63 ;
		RECT	1.57 34.485 1.62 34.615 ;
		RECT	3.02 34.46 3.15 34.64 ;
		RECT	4.87 34.485 4.92 34.615 ;
		RECT	5.9 34.485 5.95 34.615 ;
		RECT	12.79 34.485 12.84 34.615 ;
		RECT	14.29 34.46 14.42 34.64 ;
		RECT	2.18 36.455 2.23 36.585 ;
		RECT	8.56 36.455 8.61 36.585 ;
		RECT	2.18 37.435 2.23 37.565 ;
		RECT	8.56 37.435 8.61 37.565 ;
		RECT	2.18 38.42 2.23 38.55 ;
		RECT	8.56 38.42 8.61 38.55 ;
		RECT	2.18 40.39 2.23 40.52 ;
		RECT	8.56 40.39 8.61 40.52 ;
		RECT	2.18 41.37 2.23 41.5 ;
		RECT	8.56 41.37 8.61 41.5 ;
		RECT	2.18 42.355 2.23 42.485 ;
		RECT	8.56 42.355 8.61 42.485 ;
		RECT	2.18 44.33 2.23 44.46 ;
		RECT	8.56 44.33 8.61 44.46 ;
		RECT	2.18 45.31 2.23 45.44 ;
		RECT	8.56 45.31 8.61 45.44 ;
		RECT	2.18 48.26 2.23 48.39 ;
		RECT	8.56 48.26 8.61 48.39 ;
		RECT	2.18 49.735 2.23 49.865 ;
		RECT	8.56 49.735 8.61 49.865 ;
		RECT	2.18 52.685 2.23 52.815 ;
		RECT	8.56 52.685 8.61 52.815 ;
		RECT	2.18 53.675 2.23 53.805 ;
		RECT	8.56 53.675 8.61 53.805 ;
		RECT	2.18 55.64 2.23 55.77 ;
		RECT	8.56 55.64 8.61 55.77 ;
		RECT	2.18 56.625 2.23 56.755 ;
		RECT	8.56 56.625 8.61 56.755 ;
		RECT	2.18 57.61 2.23 57.74 ;
		RECT	8.56 57.61 8.61 57.74 ;
		RECT	2.18 59.575 2.23 59.705 ;
		RECT	8.56 59.575 8.61 59.705 ;
		RECT	2.18 60.56 2.23 60.69 ;
		RECT	8.56 60.56 8.61 60.69 ;
		RECT	2.18 61.545 2.23 61.675 ;
		RECT	8.56 61.545 8.61 61.675 ;
		RECT	1.57 63.515 1.62 63.645 ;
		RECT	3.02 63.49 3.15 63.67 ;
		RECT	4.87 63.515 4.92 63.645 ;
		RECT	6.375 63.515 6.425 63.645 ;
		RECT	12.79 63.515 12.84 63.645 ;
		RECT	14.29 63.49 14.42 63.67 ;
		RECT	2.18 64.495 2.23 64.625 ;
		RECT	8.56 64.495 8.61 64.625 ;
		RECT	10.27 64.495 10.32 64.625 ;
		RECT	2.18 65.48 2.23 65.61 ;
		RECT	8.56 65.48 8.61 65.61 ;
		RECT	10.27 65.48 10.32 65.61 ;
		RECT	2.18 67.45 2.23 67.58 ;
		RECT	8.56 67.45 8.61 67.58 ;
		RECT	10.27 67.45 10.32 67.58 ;
		RECT	2.18 68.435 2.23 68.565 ;
		RECT	8.56 68.435 8.61 68.565 ;
		RECT	10.27 68.435 10.32 68.565 ;
		RECT	3.06 69.455 3.11 69.585 ;
		RECT	4.87 69.455 4.92 69.585 ;
		RECT	6.375 69.455 6.425 69.585 ;
		RECT	8.975 69.455 9.025 69.585 ;
		RECT	12.79 69.455 12.84 69.585 ;
		RECT	14.33 69.455 14.38 69.585 ;
		RECT	51.115 0.425 51.295 0.555 ;
		RECT	14.965 0.655 15.015 0.785 ;
		RECT	49.725 0.655 49.775 0.785 ;
		RECT	14.765 0.655 14.815 0.785 ;
		RECT	49.925 0.655 49.975 0.785 ;
		RECT	50.94 0.425 50.99 0.555 ;
		RECT	51.115 100.385 51.295 100.515 ;
		RECT	14.965 100.155 15.015 100.285 ;
		RECT	49.725 100.155 49.775 100.285 ;
		RECT	14.765 100.155 14.815 100.285 ;
		RECT	49.925 100.155 49.975 100.285 ;
		RECT	50.94 100.385 50.99 100.515 ;
		RECT	14.565 3.305 14.615 3.435 ;
		RECT	50.125 3.305 50.175 3.435 ;
		RECT	14.765 3.535 14.815 3.665 ;
		RECT	14.765 1.115 14.815 1.245 ;
		RECT	49.925 3.535 49.975 3.665 ;
		RECT	49.925 1.115 49.975 1.245 ;
		RECT	14.965 3.535 15.015 3.665 ;
		RECT	14.965 1.115 15.015 1.245 ;
		RECT	49.725 3.535 49.775 3.665 ;
		RECT	49.725 1.115 49.775 1.245 ;
		RECT	14.565 26.345 14.615 26.475 ;
		RECT	50.125 26.345 50.175 26.475 ;
		RECT	14.765 26.575 14.815 26.705 ;
		RECT	14.765 24.155 14.815 24.285 ;
		RECT	49.925 26.575 49.975 26.705 ;
		RECT	49.925 24.155 49.975 24.285 ;
		RECT	14.965 26.575 15.015 26.705 ;
		RECT	14.965 24.155 15.015 24.285 ;
		RECT	49.725 26.575 49.775 26.705 ;
		RECT	49.725 24.155 49.775 24.285 ;
		RECT	14.565 23.465 14.615 23.595 ;
		RECT	50.125 23.465 50.175 23.595 ;
		RECT	14.765 23.695 14.815 23.825 ;
		RECT	14.765 21.275 14.815 21.405 ;
		RECT	49.925 23.695 49.975 23.825 ;
		RECT	49.925 21.275 49.975 21.405 ;
		RECT	14.965 23.695 15.015 23.825 ;
		RECT	14.965 21.275 15.015 21.405 ;
		RECT	49.725 23.695 49.775 23.825 ;
		RECT	49.725 21.275 49.775 21.405 ;
		RECT	14.565 20.585 14.615 20.715 ;
		RECT	50.125 20.585 50.175 20.715 ;
		RECT	14.765 20.815 14.815 20.945 ;
		RECT	14.765 18.395 14.815 18.525 ;
		RECT	49.925 20.815 49.975 20.945 ;
		RECT	49.925 18.395 49.975 18.525 ;
		RECT	14.965 20.815 15.015 20.945 ;
		RECT	14.965 18.395 15.015 18.525 ;
		RECT	49.725 20.815 49.775 20.945 ;
		RECT	49.725 18.395 49.775 18.525 ;
		RECT	14.565 17.705 14.615 17.835 ;
		RECT	50.125 17.705 50.175 17.835 ;
		RECT	14.765 17.935 14.815 18.065 ;
		RECT	14.765 15.515 14.815 15.645 ;
		RECT	49.925 17.935 49.975 18.065 ;
		RECT	49.925 15.515 49.975 15.645 ;
		RECT	14.965 17.935 15.015 18.065 ;
		RECT	14.965 15.515 15.015 15.645 ;
		RECT	49.725 17.935 49.775 18.065 ;
		RECT	49.725 15.515 49.775 15.645 ;
		RECT	14.565 14.825 14.615 14.955 ;
		RECT	50.125 14.825 50.175 14.955 ;
		RECT	14.765 15.055 14.815 15.185 ;
		RECT	14.765 12.635 14.815 12.765 ;
		RECT	49.925 15.055 49.975 15.185 ;
		RECT	49.925 12.635 49.975 12.765 ;
		RECT	14.965 15.055 15.015 15.185 ;
		RECT	14.965 12.635 15.015 12.765 ;
		RECT	49.725 15.055 49.775 15.185 ;
		RECT	49.725 12.635 49.775 12.765 ;
		RECT	14.565 11.945 14.615 12.075 ;
		RECT	50.125 11.945 50.175 12.075 ;
		RECT	14.765 12.175 14.815 12.305 ;
		RECT	14.765 9.755 14.815 9.885 ;
		RECT	49.925 12.175 49.975 12.305 ;
		RECT	49.925 9.755 49.975 9.885 ;
		RECT	14.965 12.175 15.015 12.305 ;
		RECT	14.965 9.755 15.015 9.885 ;
		RECT	49.725 12.175 49.775 12.305 ;
		RECT	49.725 9.755 49.775 9.885 ;
		RECT	14.565 9.065 14.615 9.195 ;
		RECT	50.125 9.065 50.175 9.195 ;
		RECT	14.765 9.295 14.815 9.425 ;
		RECT	14.765 6.875 14.815 7.005 ;
		RECT	49.925 9.295 49.975 9.425 ;
		RECT	49.925 6.875 49.975 7.005 ;
		RECT	14.965 9.295 15.015 9.425 ;
		RECT	14.965 6.875 15.015 7.005 ;
		RECT	49.725 9.295 49.775 9.425 ;
		RECT	49.725 6.875 49.775 7.005 ;
		RECT	14.565 6.185 14.615 6.315 ;
		RECT	50.125 6.185 50.175 6.315 ;
		RECT	14.765 6.415 14.815 6.545 ;
		RECT	14.765 3.995 14.815 4.125 ;
		RECT	49.925 6.415 49.975 6.545 ;
		RECT	49.925 3.995 49.975 4.125 ;
		RECT	14.965 6.415 15.015 6.545 ;
		RECT	14.965 3.995 15.015 4.125 ;
		RECT	49.725 6.415 49.775 6.545 ;
		RECT	49.725 3.995 49.775 4.125 ;
		RECT	50.325 23.695 50.505 23.825 ;
		RECT	51.115 23.465 51.295 23.595 ;
		RECT	50.325 21.275 50.505 21.405 ;
		RECT	50.67 21.045 50.72 21.175 ;
		RECT	50.325 20.815 50.505 20.945 ;
		RECT	51.115 20.585 51.295 20.715 ;
		RECT	50.325 18.395 50.505 18.525 ;
		RECT	50.67 18.165 50.72 18.295 ;
		RECT	50.325 17.935 50.505 18.065 ;
		RECT	51.115 17.705 51.295 17.835 ;
		RECT	50.325 15.515 50.505 15.645 ;
		RECT	50.67 15.285 50.72 15.415 ;
		RECT	50.325 15.055 50.505 15.185 ;
		RECT	51.115 14.825 51.295 14.955 ;
		RECT	50.325 12.635 50.505 12.765 ;
		RECT	50.67 12.405 50.72 12.535 ;
		RECT	50.325 12.175 50.505 12.305 ;
		RECT	51.115 11.945 51.295 12.075 ;
		RECT	50.325 9.755 50.505 9.885 ;
		RECT	50.67 9.525 50.72 9.655 ;
		RECT	50.325 9.295 50.505 9.425 ;
		RECT	51.115 9.065 51.295 9.195 ;
		RECT	50.325 6.875 50.505 7.005 ;
		RECT	50.67 6.645 50.72 6.775 ;
		RECT	50.325 6.415 50.505 6.545 ;
		RECT	51.115 6.185 51.295 6.315 ;
		RECT	50.325 3.995 50.505 4.125 ;
		RECT	50.67 3.765 50.72 3.895 ;
		RECT	50.325 3.535 50.505 3.665 ;
		RECT	51.115 3.305 51.295 3.435 ;
		RECT	50.325 1.115 50.505 1.245 ;
		RECT	50.67 0.885 50.72 1.015 ;
		RECT	50.325 26.575 50.505 26.705 ;
		RECT	51.115 26.345 51.295 26.475 ;
		RECT	50.325 24.155 50.505 24.285 ;
		RECT	50.67 23.925 50.72 24.055 ;
		RECT	14.565 97.505 14.615 97.635 ;
		RECT	50.125 97.505 50.175 97.635 ;
		RECT	14.765 97.275 14.815 97.405 ;
		RECT	14.765 99.695 14.815 99.825 ;
		RECT	49.925 97.275 49.975 97.405 ;
		RECT	49.925 99.695 49.975 99.825 ;
		RECT	14.965 97.275 15.015 97.405 ;
		RECT	14.965 99.695 15.015 99.825 ;
		RECT	49.725 97.275 49.775 97.405 ;
		RECT	49.725 99.695 49.775 99.825 ;
		RECT	14.565 71.585 14.615 71.715 ;
		RECT	50.125 71.585 50.175 71.715 ;
		RECT	14.765 71.355 14.815 71.485 ;
		RECT	14.765 73.775 14.815 73.905 ;
		RECT	49.925 71.355 49.975 71.485 ;
		RECT	49.925 73.775 49.975 73.905 ;
		RECT	14.965 71.355 15.015 71.485 ;
		RECT	14.965 73.775 15.015 73.905 ;
		RECT	49.725 71.355 49.775 71.485 ;
		RECT	49.725 73.775 49.775 73.905 ;
		RECT	14.565 74.465 14.615 74.595 ;
		RECT	50.125 74.465 50.175 74.595 ;
		RECT	14.765 74.235 14.815 74.365 ;
		RECT	14.765 76.655 14.815 76.785 ;
		RECT	49.925 74.235 49.975 74.365 ;
		RECT	49.925 76.655 49.975 76.785 ;
		RECT	14.965 74.235 15.015 74.365 ;
		RECT	14.965 76.655 15.015 76.785 ;
		RECT	49.725 74.235 49.775 74.365 ;
		RECT	49.725 76.655 49.775 76.785 ;
		RECT	14.565 77.345 14.615 77.475 ;
		RECT	50.125 77.345 50.175 77.475 ;
		RECT	14.765 77.115 14.815 77.245 ;
		RECT	14.765 79.535 14.815 79.665 ;
		RECT	49.925 77.115 49.975 77.245 ;
		RECT	49.925 79.535 49.975 79.665 ;
		RECT	14.965 77.115 15.015 77.245 ;
		RECT	14.965 79.535 15.015 79.665 ;
		RECT	49.725 77.115 49.775 77.245 ;
		RECT	49.725 79.535 49.775 79.665 ;
		RECT	14.565 80.225 14.615 80.355 ;
		RECT	50.125 80.225 50.175 80.355 ;
		RECT	14.765 79.995 14.815 80.125 ;
		RECT	14.765 82.415 14.815 82.545 ;
		RECT	49.925 79.995 49.975 80.125 ;
		RECT	49.925 82.415 49.975 82.545 ;
		RECT	14.965 79.995 15.015 80.125 ;
		RECT	14.965 82.415 15.015 82.545 ;
		RECT	49.725 79.995 49.775 80.125 ;
		RECT	49.725 82.415 49.775 82.545 ;
		RECT	14.565 83.105 14.615 83.235 ;
		RECT	50.125 83.105 50.175 83.235 ;
		RECT	14.765 82.875 14.815 83.005 ;
		RECT	14.765 85.295 14.815 85.425 ;
		RECT	49.925 82.875 49.975 83.005 ;
		RECT	49.925 85.295 49.975 85.425 ;
		RECT	14.965 82.875 15.015 83.005 ;
		RECT	14.965 85.295 15.015 85.425 ;
		RECT	49.725 82.875 49.775 83.005 ;
		RECT	49.725 85.295 49.775 85.425 ;
		RECT	14.565 85.985 14.615 86.115 ;
		RECT	50.125 85.985 50.175 86.115 ;
		RECT	14.765 85.755 14.815 85.885 ;
		RECT	14.765 88.175 14.815 88.305 ;
		RECT	49.925 85.755 49.975 85.885 ;
		RECT	49.925 88.175 49.975 88.305 ;
		RECT	14.965 85.755 15.015 85.885 ;
		RECT	14.965 88.175 15.015 88.305 ;
		RECT	49.725 85.755 49.775 85.885 ;
		RECT	49.725 88.175 49.775 88.305 ;
		RECT	14.565 88.865 14.615 88.995 ;
		RECT	50.125 88.865 50.175 88.995 ;
		RECT	14.765 88.635 14.815 88.765 ;
		RECT	14.765 91.055 14.815 91.185 ;
		RECT	49.925 88.635 49.975 88.765 ;
		RECT	49.925 91.055 49.975 91.185 ;
		RECT	14.965 88.635 15.015 88.765 ;
		RECT	14.965 91.055 15.015 91.185 ;
		RECT	49.725 88.635 49.775 88.765 ;
		RECT	49.725 91.055 49.775 91.185 ;
		RECT	14.565 91.745 14.615 91.875 ;
		RECT	50.125 91.745 50.175 91.875 ;
		RECT	14.765 91.515 14.815 91.645 ;
		RECT	14.765 93.935 14.815 94.065 ;
		RECT	49.925 91.515 49.975 91.645 ;
		RECT	49.925 93.935 49.975 94.065 ;
		RECT	14.965 91.515 15.015 91.645 ;
		RECT	14.965 93.935 15.015 94.065 ;
		RECT	49.725 91.515 49.775 91.645 ;
		RECT	49.725 93.935 49.775 94.065 ;
		RECT	14.565 94.625 14.615 94.755 ;
		RECT	50.125 94.625 50.175 94.755 ;
		RECT	14.765 94.395 14.815 94.525 ;
		RECT	14.765 96.815 14.815 96.945 ;
		RECT	49.925 94.395 49.975 94.525 ;
		RECT	49.925 96.815 49.975 96.945 ;
		RECT	14.965 94.395 15.015 94.525 ;
		RECT	14.965 96.815 15.015 96.945 ;
		RECT	49.725 94.395 49.775 94.525 ;
		RECT	49.725 96.815 49.775 96.945 ;
		RECT	50.325 74.235 50.505 74.365 ;
		RECT	51.115 74.465 51.295 74.595 ;
		RECT	50.325 76.655 50.505 76.785 ;
		RECT	50.67 76.885 50.72 77.015 ;
		RECT	50.325 77.115 50.505 77.245 ;
		RECT	51.115 77.345 51.295 77.475 ;
		RECT	50.325 79.535 50.505 79.665 ;
		RECT	50.67 79.765 50.72 79.895 ;
		RECT	50.325 79.995 50.505 80.125 ;
		RECT	51.115 80.225 51.295 80.355 ;
		RECT	50.325 82.415 50.505 82.545 ;
		RECT	50.67 82.645 50.72 82.775 ;
		RECT	50.325 82.875 50.505 83.005 ;
		RECT	51.115 83.105 51.295 83.235 ;
		RECT	50.325 85.295 50.505 85.425 ;
		RECT	50.67 85.525 50.72 85.655 ;
		RECT	50.325 85.755 50.505 85.885 ;
		RECT	51.115 85.985 51.295 86.115 ;
		RECT	50.325 88.175 50.505 88.305 ;
		RECT	50.67 88.405 50.72 88.535 ;
		RECT	50.325 88.635 50.505 88.765 ;
		RECT	51.115 88.865 51.295 88.995 ;
		RECT	50.325 91.055 50.505 91.185 ;
		RECT	50.67 91.285 50.72 91.415 ;
		RECT	50.325 91.515 50.505 91.645 ;
		RECT	51.115 91.745 51.295 91.875 ;
		RECT	50.325 93.935 50.505 94.065 ;
		RECT	50.67 94.165 50.72 94.295 ;
		RECT	50.325 94.395 50.505 94.525 ;
		RECT	51.115 94.625 51.295 94.755 ;
		RECT	50.325 96.815 50.505 96.945 ;
		RECT	50.67 97.045 50.72 97.175 ;
		RECT	50.325 97.275 50.505 97.405 ;
		RECT	51.115 97.505 51.295 97.635 ;
		RECT	50.325 99.695 50.505 99.825 ;
		RECT	50.67 99.925 50.72 100.055 ;
		RECT	50.325 71.355 50.505 71.485 ;
		RECT	51.115 71.585 51.295 71.715 ;
		RECT	50.325 73.775 50.505 73.905 ;
		RECT	50.67 74.005 50.72 74.135 ;
		RECT	6.22 20.815 6.27 20.945 ;
		RECT	7.5 20.815 7.55 20.945 ;
		RECT	9.04 20.815 9.09 20.945 ;
		RECT	9.315 20.815 9.365 20.945 ;
		RECT	9.72 20.815 9.77 20.945 ;
		RECT	11.025 20.815 11.075 20.945 ;
		RECT	12.79 20.815 12.84 20.945 ;
		RECT	6.225 18.395 6.275 18.525 ;
		RECT	7.5 18.395 7.55 18.525 ;
		RECT	9.04 18.395 9.09 18.525 ;
		RECT	9.315 18.395 9.365 18.525 ;
		RECT	11.025 18.395 11.075 18.525 ;
		RECT	12.79 18.395 12.84 18.525 ;
		RECT	7.18 18.165 7.23 18.295 ;
		RECT	14.14 18.165 14.19 18.295 ;
		RECT	8.56 20.815 8.61 20.945 ;
		RECT	10.27 20.815 10.32 20.945 ;
		RECT	8.56 18.395 8.61 18.525 ;
		RECT	10.27 18.395 10.32 18.525 ;
		RECT	6.22 17.935 6.27 18.065 ;
		RECT	7.5 17.935 7.55 18.065 ;
		RECT	9.04 17.935 9.09 18.065 ;
		RECT	9.315 17.935 9.365 18.065 ;
		RECT	9.72 17.935 9.77 18.065 ;
		RECT	11.025 17.935 11.075 18.065 ;
		RECT	12.79 17.935 12.84 18.065 ;
		RECT	6.225 15.515 6.275 15.645 ;
		RECT	7.5 15.515 7.55 15.645 ;
		RECT	9.04 15.515 9.09 15.645 ;
		RECT	9.315 15.515 9.365 15.645 ;
		RECT	11.025 15.515 11.075 15.645 ;
		RECT	12.79 15.515 12.84 15.645 ;
		RECT	7.18 15.285 7.23 15.415 ;
		RECT	14.14 15.285 14.19 15.415 ;
		RECT	8.56 17.935 8.61 18.065 ;
		RECT	10.27 17.935 10.32 18.065 ;
		RECT	8.56 15.515 8.61 15.645 ;
		RECT	10.27 15.515 10.32 15.645 ;
		RECT	6.22 15.055 6.27 15.185 ;
		RECT	7.5 15.055 7.55 15.185 ;
		RECT	9.04 15.055 9.09 15.185 ;
		RECT	9.315 15.055 9.365 15.185 ;
		RECT	9.72 15.055 9.77 15.185 ;
		RECT	11.025 15.055 11.075 15.185 ;
		RECT	12.79 15.055 12.84 15.185 ;
		RECT	6.225 12.635 6.275 12.765 ;
		RECT	7.5 12.635 7.55 12.765 ;
		RECT	9.04 12.635 9.09 12.765 ;
		RECT	9.315 12.635 9.365 12.765 ;
		RECT	11.025 12.635 11.075 12.765 ;
		RECT	12.79 12.635 12.84 12.765 ;
		RECT	7.18 12.405 7.23 12.535 ;
		RECT	14.14 12.405 14.19 12.535 ;
		RECT	8.56 15.055 8.61 15.185 ;
		RECT	10.27 15.055 10.32 15.185 ;
		RECT	8.56 12.635 8.61 12.765 ;
		RECT	10.27 12.635 10.32 12.765 ;
		RECT	6.22 12.175 6.27 12.305 ;
		RECT	7.5 12.175 7.55 12.305 ;
		RECT	9.04 12.175 9.09 12.305 ;
		RECT	9.315 12.175 9.365 12.305 ;
		RECT	9.72 12.175 9.77 12.305 ;
		RECT	11.025 12.175 11.075 12.305 ;
		RECT	12.79 12.175 12.84 12.305 ;
		RECT	6.225 9.755 6.275 9.885 ;
		RECT	7.5 9.755 7.55 9.885 ;
		RECT	9.04 9.755 9.09 9.885 ;
		RECT	9.315 9.755 9.365 9.885 ;
		RECT	11.025 9.755 11.075 9.885 ;
		RECT	12.79 9.755 12.84 9.885 ;
		RECT	7.18 9.525 7.23 9.655 ;
		RECT	14.14 9.525 14.19 9.655 ;
		RECT	8.56 12.175 8.61 12.305 ;
		RECT	10.27 12.175 10.32 12.305 ;
		RECT	8.56 9.755 8.61 9.885 ;
		RECT	10.27 9.755 10.32 9.885 ;
		RECT	6.22 9.295 6.27 9.425 ;
		RECT	7.5 9.295 7.55 9.425 ;
		RECT	9.04 9.295 9.09 9.425 ;
		RECT	9.315 9.295 9.365 9.425 ;
		RECT	9.72 9.295 9.77 9.425 ;
		RECT	11.025 9.295 11.075 9.425 ;
		RECT	12.79 9.295 12.84 9.425 ;
		RECT	6.225 6.875 6.275 7.005 ;
		RECT	7.5 6.875 7.55 7.005 ;
		RECT	9.04 6.875 9.09 7.005 ;
		RECT	9.315 6.875 9.365 7.005 ;
		RECT	11.025 6.875 11.075 7.005 ;
		RECT	12.79 6.875 12.84 7.005 ;
		RECT	7.18 6.645 7.23 6.775 ;
		RECT	14.14 6.645 14.19 6.775 ;
		RECT	8.56 9.295 8.61 9.425 ;
		RECT	10.27 9.295 10.32 9.425 ;
		RECT	8.56 6.875 8.61 7.005 ;
		RECT	10.27 6.875 10.32 7.005 ;
		RECT	6.22 6.415 6.27 6.545 ;
		RECT	7.5 6.415 7.55 6.545 ;
		RECT	9.04 6.415 9.09 6.545 ;
		RECT	9.315 6.415 9.365 6.545 ;
		RECT	9.72 6.415 9.77 6.545 ;
		RECT	11.025 6.415 11.075 6.545 ;
		RECT	12.79 6.415 12.84 6.545 ;
		RECT	6.225 3.995 6.275 4.125 ;
		RECT	7.5 3.995 7.55 4.125 ;
		RECT	9.04 3.995 9.09 4.125 ;
		RECT	9.315 3.995 9.365 4.125 ;
		RECT	11.025 3.995 11.075 4.125 ;
		RECT	12.79 3.995 12.84 4.125 ;
		RECT	7.18 3.765 7.23 3.895 ;
		RECT	14.14 3.765 14.19 3.895 ;
		RECT	8.56 6.415 8.61 6.545 ;
		RECT	10.27 6.415 10.32 6.545 ;
		RECT	8.56 3.995 8.61 4.125 ;
		RECT	10.27 3.995 10.32 4.125 ;
		RECT	6.22 3.535 6.27 3.665 ;
		RECT	7.5 3.535 7.55 3.665 ;
		RECT	9.04 3.535 9.09 3.665 ;
		RECT	9.315 3.535 9.365 3.665 ;
		RECT	9.72 3.535 9.77 3.665 ;
		RECT	11.025 3.535 11.075 3.665 ;
		RECT	12.79 3.535 12.84 3.665 ;
		RECT	6.225 1.115 6.275 1.245 ;
		RECT	7.5 1.115 7.55 1.245 ;
		RECT	9.04 1.115 9.09 1.245 ;
		RECT	9.315 1.115 9.365 1.245 ;
		RECT	11.025 1.115 11.075 1.245 ;
		RECT	12.79 1.115 12.84 1.245 ;
		RECT	7.18 0.885 7.23 1.015 ;
		RECT	14.14 0.885 14.19 1.015 ;
		RECT	8.56 3.535 8.61 3.665 ;
		RECT	10.27 3.535 10.32 3.665 ;
		RECT	8.56 1.115 8.61 1.245 ;
		RECT	10.27 1.115 10.32 1.245 ;
		RECT	6.22 26.575 6.27 26.705 ;
		RECT	7.5 26.575 7.55 26.705 ;
		RECT	9.04 26.575 9.09 26.705 ;
		RECT	9.315 26.575 9.365 26.705 ;
		RECT	9.72 26.575 9.77 26.705 ;
		RECT	11.025 26.575 11.075 26.705 ;
		RECT	12.79 26.575 12.84 26.705 ;
		RECT	6.225 24.155 6.275 24.285 ;
		RECT	7.5 24.155 7.55 24.285 ;
		RECT	9.04 24.155 9.09 24.285 ;
		RECT	9.315 24.155 9.365 24.285 ;
		RECT	11.025 24.155 11.075 24.285 ;
		RECT	12.79 24.155 12.84 24.285 ;
		RECT	7.18 23.925 7.23 24.055 ;
		RECT	14.14 23.925 14.19 24.055 ;
		RECT	8.56 26.575 8.61 26.705 ;
		RECT	10.27 26.575 10.32 26.705 ;
		RECT	8.56 24.155 8.61 24.285 ;
		RECT	10.27 24.155 10.32 24.285 ;
		RECT	6.22 23.695 6.27 23.825 ;
		RECT	7.5 23.695 7.55 23.825 ;
		RECT	9.04 23.695 9.09 23.825 ;
		RECT	9.315 23.695 9.365 23.825 ;
		RECT	9.72 23.695 9.77 23.825 ;
		RECT	11.025 23.695 11.075 23.825 ;
		RECT	12.79 23.695 12.84 23.825 ;
		RECT	6.225 21.275 6.275 21.405 ;
		RECT	7.5 21.275 7.55 21.405 ;
		RECT	9.04 21.275 9.09 21.405 ;
		RECT	9.315 21.275 9.365 21.405 ;
		RECT	11.025 21.275 11.075 21.405 ;
		RECT	12.79 21.275 12.84 21.405 ;
		RECT	7.18 21.045 7.23 21.175 ;
		RECT	14.14 21.045 14.19 21.175 ;
		RECT	8.56 23.695 8.61 23.825 ;
		RECT	10.27 23.695 10.32 23.825 ;
		RECT	8.56 21.275 8.61 21.405 ;
		RECT	10.27 21.275 10.32 21.405 ;
		RECT	14.33 23.695 14.38 23.825 ;
		RECT	6.22 23.235 6.27 23.365 ;
		RECT	7.5 23.235 7.55 23.365 ;
		RECT	9.04 23.235 9.09 23.365 ;
		RECT	9.315 23.235 9.365 23.365 ;
		RECT	9.72 23.235 9.77 23.365 ;
		RECT	11.025 23.235 11.075 23.365 ;
		RECT	12.79 23.235 12.84 23.365 ;
		RECT	14.33 21.275 14.38 21.405 ;
		RECT	5.675 21.045 5.725 21.175 ;
		RECT	6.065 21.045 6.115 21.175 ;
		RECT	6.725 21.045 6.775 21.175 ;
		RECT	8.42 21.045 8.47 21.175 ;
		RECT	8.77 21.045 8.82 21.175 ;
		RECT	11.555 21.045 11.605 21.175 ;
		RECT	11.815 21.045 11.865 21.175 ;
		RECT	12.52 21.045 12.57 21.175 ;
		RECT	13.98 21.045 14.03 21.175 ;
		RECT	14.33 20.815 14.38 20.945 ;
		RECT	6.22 20.355 6.27 20.485 ;
		RECT	7.5 20.355 7.55 20.485 ;
		RECT	9.04 20.355 9.09 20.485 ;
		RECT	9.315 20.355 9.365 20.485 ;
		RECT	9.72 20.355 9.77 20.485 ;
		RECT	11.025 20.355 11.075 20.485 ;
		RECT	12.79 20.355 12.84 20.485 ;
		RECT	14.33 18.395 14.38 18.525 ;
		RECT	5.675 18.165 5.725 18.295 ;
		RECT	6.065 18.165 6.115 18.295 ;
		RECT	6.725 18.165 6.775 18.295 ;
		RECT	8.42 18.165 8.47 18.295 ;
		RECT	8.77 18.165 8.82 18.295 ;
		RECT	11.555 18.165 11.605 18.295 ;
		RECT	11.815 18.165 11.865 18.295 ;
		RECT	12.52 18.165 12.57 18.295 ;
		RECT	13.98 18.165 14.03 18.295 ;
		RECT	14.33 17.935 14.38 18.065 ;
		RECT	6.22 17.475 6.27 17.605 ;
		RECT	7.5 17.475 7.55 17.605 ;
		RECT	9.04 17.475 9.09 17.605 ;
		RECT	9.315 17.475 9.365 17.605 ;
		RECT	9.72 17.475 9.77 17.605 ;
		RECT	11.025 17.475 11.075 17.605 ;
		RECT	12.79 17.475 12.84 17.605 ;
		RECT	14.33 15.515 14.38 15.645 ;
		RECT	5.675 15.285 5.725 15.415 ;
		RECT	6.065 15.285 6.115 15.415 ;
		RECT	6.725 15.285 6.775 15.415 ;
		RECT	8.42 15.285 8.47 15.415 ;
		RECT	8.77 15.285 8.82 15.415 ;
		RECT	11.555 15.285 11.605 15.415 ;
		RECT	11.815 15.285 11.865 15.415 ;
		RECT	12.52 15.285 12.57 15.415 ;
		RECT	13.98 15.285 14.03 15.415 ;
		RECT	14.33 15.055 14.38 15.185 ;
		RECT	6.22 14.595 6.27 14.725 ;
		RECT	7.5 14.595 7.55 14.725 ;
		RECT	9.04 14.595 9.09 14.725 ;
		RECT	9.315 14.595 9.365 14.725 ;
		RECT	9.72 14.595 9.77 14.725 ;
		RECT	11.025 14.595 11.075 14.725 ;
		RECT	12.79 14.595 12.84 14.725 ;
		RECT	14.33 12.635 14.38 12.765 ;
		RECT	5.675 12.405 5.725 12.535 ;
		RECT	6.065 12.405 6.115 12.535 ;
		RECT	6.725 12.405 6.775 12.535 ;
		RECT	8.42 12.405 8.47 12.535 ;
		RECT	8.77 12.405 8.82 12.535 ;
		RECT	11.555 12.405 11.605 12.535 ;
		RECT	11.815 12.405 11.865 12.535 ;
		RECT	12.52 12.405 12.57 12.535 ;
		RECT	13.98 12.405 14.03 12.535 ;
		RECT	14.33 12.175 14.38 12.305 ;
		RECT	6.22 11.715 6.27 11.845 ;
		RECT	7.5 11.715 7.55 11.845 ;
		RECT	9.04 11.715 9.09 11.845 ;
		RECT	9.315 11.715 9.365 11.845 ;
		RECT	9.72 11.715 9.77 11.845 ;
		RECT	11.025 11.715 11.075 11.845 ;
		RECT	12.79 11.715 12.84 11.845 ;
		RECT	14.33 9.755 14.38 9.885 ;
		RECT	5.675 9.525 5.725 9.655 ;
		RECT	6.065 9.525 6.115 9.655 ;
		RECT	6.725 9.525 6.775 9.655 ;
		RECT	8.42 9.525 8.47 9.655 ;
		RECT	8.77 9.525 8.82 9.655 ;
		RECT	11.555 9.525 11.605 9.655 ;
		RECT	11.815 9.525 11.865 9.655 ;
		RECT	12.52 9.525 12.57 9.655 ;
		RECT	13.98 9.525 14.03 9.655 ;
		RECT	14.33 9.295 14.38 9.425 ;
		RECT	6.22 8.835 6.27 8.965 ;
		RECT	7.5 8.835 7.55 8.965 ;
		RECT	9.04 8.835 9.09 8.965 ;
		RECT	9.315 8.835 9.365 8.965 ;
		RECT	9.72 8.835 9.77 8.965 ;
		RECT	11.025 8.835 11.075 8.965 ;
		RECT	12.79 8.835 12.84 8.965 ;
		RECT	14.33 6.875 14.38 7.005 ;
		RECT	5.675 6.645 5.725 6.775 ;
		RECT	6.065 6.645 6.115 6.775 ;
		RECT	6.725 6.645 6.775 6.775 ;
		RECT	8.42 6.645 8.47 6.775 ;
		RECT	8.77 6.645 8.82 6.775 ;
		RECT	11.555 6.645 11.605 6.775 ;
		RECT	11.815 6.645 11.865 6.775 ;
		RECT	12.52 6.645 12.57 6.775 ;
		RECT	13.98 6.645 14.03 6.775 ;
		RECT	14.33 6.415 14.38 6.545 ;
		RECT	6.22 5.955 6.27 6.085 ;
		RECT	7.5 5.955 7.55 6.085 ;
		RECT	9.04 5.955 9.09 6.085 ;
		RECT	9.315 5.955 9.365 6.085 ;
		RECT	9.72 5.955 9.77 6.085 ;
		RECT	11.025 5.955 11.075 6.085 ;
		RECT	12.79 5.955 12.84 6.085 ;
		RECT	14.33 3.995 14.38 4.125 ;
		RECT	5.675 3.765 5.725 3.895 ;
		RECT	6.065 3.765 6.115 3.895 ;
		RECT	6.725 3.765 6.775 3.895 ;
		RECT	8.42 3.765 8.47 3.895 ;
		RECT	8.77 3.765 8.82 3.895 ;
		RECT	11.555 3.765 11.605 3.895 ;
		RECT	11.815 3.765 11.865 3.895 ;
		RECT	12.52 3.765 12.57 3.895 ;
		RECT	13.98 3.765 14.03 3.895 ;
		RECT	14.33 3.535 14.38 3.665 ;
		RECT	6.22 3.075 6.27 3.205 ;
		RECT	7.5 3.075 7.55 3.205 ;
		RECT	9.04 3.075 9.09 3.205 ;
		RECT	9.315 3.075 9.365 3.205 ;
		RECT	9.72 3.075 9.77 3.205 ;
		RECT	11.025 3.075 11.075 3.205 ;
		RECT	12.79 3.075 12.84 3.205 ;
		RECT	14.33 1.115 14.38 1.245 ;
		RECT	5.675 0.885 5.725 1.015 ;
		RECT	6.065 0.885 6.115 1.015 ;
		RECT	6.725 0.885 6.775 1.015 ;
		RECT	8.42 0.885 8.47 1.015 ;
		RECT	8.77 0.885 8.82 1.015 ;
		RECT	11.555 0.885 11.605 1.015 ;
		RECT	11.815 0.885 11.865 1.015 ;
		RECT	12.52 0.885 12.57 1.015 ;
		RECT	13.98 0.885 14.03 1.015 ;
		RECT	14.33 26.575 14.38 26.705 ;
		RECT	6.22 26.115 6.27 26.245 ;
		RECT	7.5 26.115 7.55 26.245 ;
		RECT	9.04 26.115 9.09 26.245 ;
		RECT	9.315 26.115 9.365 26.245 ;
		RECT	9.72 26.115 9.77 26.245 ;
		RECT	11.025 26.115 11.075 26.245 ;
		RECT	12.79 26.115 12.84 26.245 ;
		RECT	14.33 24.155 14.38 24.285 ;
		RECT	5.675 23.925 5.725 24.055 ;
		RECT	6.065 23.925 6.115 24.055 ;
		RECT	6.725 23.925 6.775 24.055 ;
		RECT	8.42 23.925 8.47 24.055 ;
		RECT	8.77 23.925 8.82 24.055 ;
		RECT	11.555 23.925 11.605 24.055 ;
		RECT	11.815 23.925 11.865 24.055 ;
		RECT	12.52 23.925 12.57 24.055 ;
		RECT	13.98 23.925 14.03 24.055 ;
		RECT	13.98 0.195 14.03 0.325 ;
		RECT	1.57 0.195 1.62 0.325 ;
		RECT	2.485 0.195 2.665 0.325 ;
		RECT	3.84 0.195 3.89 0.325 ;
		RECT	7.19 0.195 7.24 0.325 ;
		RECT	14.14 0.195 14.19 0.325 ;
		RECT	13.8 0.425 13.85 0.555 ;
		RECT	8.56 0.655 8.61 0.785 ;
		RECT	10.27 0.655 10.32 0.785 ;
		RECT	0.435 0.655 0.485 0.785 ;
		RECT	0.62 0.195 0.67 0.325 ;
		RECT	3.65 0.195 3.7 0.325 ;
		RECT	2.18 0.655 2.23 0.785 ;
		RECT	0.9 21.045 0.95 21.175 ;
		RECT	0.9 18.165 0.95 18.295 ;
		RECT	0.9 15.285 0.95 15.415 ;
		RECT	0.9 12.405 0.95 12.535 ;
		RECT	0.9 9.525 0.95 9.655 ;
		RECT	0.9 6.645 0.95 6.775 ;
		RECT	0.9 3.765 0.95 3.895 ;
		RECT	0.9 0.885 0.95 1.015 ;
		RECT	0.9 23.925 0.95 24.055 ;
		RECT	3.65 23.925 3.7 24.055 ;
		RECT	3.65 21.045 3.7 21.175 ;
		RECT	3.65 18.165 3.7 18.295 ;
		RECT	3.65 15.285 3.7 15.415 ;
		RECT	3.65 12.405 3.7 12.535 ;
		RECT	3.65 9.525 3.7 9.655 ;
		RECT	3.65 6.645 3.7 6.775 ;
		RECT	3.65 3.765 3.7 3.895 ;
		RECT	3.65 0.885 3.7 1.015 ;
		RECT	2.18 26.575 2.23 26.705 ;
		RECT	2.18 24.155 2.23 24.285 ;
		RECT	2.18 23.695 2.23 23.825 ;
		RECT	2.18 21.275 2.23 21.405 ;
		RECT	2.18 20.815 2.23 20.945 ;
		RECT	2.18 18.395 2.23 18.525 ;
		RECT	2.18 17.935 2.23 18.065 ;
		RECT	2.18 15.515 2.23 15.645 ;
		RECT	2.18 15.055 2.23 15.185 ;
		RECT	2.18 12.635 2.23 12.765 ;
		RECT	2.18 12.175 2.23 12.305 ;
		RECT	2.18 9.755 2.23 9.885 ;
		RECT	2.18 9.295 2.23 9.425 ;
		RECT	2.18 6.875 2.23 7.005 ;
		RECT	2.18 6.415 2.23 6.545 ;
		RECT	2.18 3.995 2.23 4.125 ;
		RECT	2.18 3.535 2.23 3.665 ;
		RECT	2.18 1.115 2.23 1.245 ;
		RECT	3.06 23.695 3.11 23.825 ;
		RECT	1.085 23.235 1.135 23.365 ;
		RECT	1.405 23.275 1.455 23.325 ;
		RECT	4.47 23.275 4.6 23.325 ;
		RECT	3.06 21.275 3.11 21.405 ;
		RECT	1.57 21.045 1.62 21.175 ;
		RECT	2.58 21.045 2.63 21.175 ;
		RECT	3.84 21.045 3.89 21.175 ;
		RECT	5.675 21.045 5.725 21.175 ;
		RECT	3.06 20.815 3.11 20.945 ;
		RECT	1.085 20.355 1.135 20.485 ;
		RECT	1.405 20.395 1.455 20.445 ;
		RECT	4.47 20.395 4.6 20.445 ;
		RECT	3.06 18.395 3.11 18.525 ;
		RECT	1.57 18.165 1.62 18.295 ;
		RECT	2.58 18.165 2.63 18.295 ;
		RECT	3.84 18.165 3.89 18.295 ;
		RECT	5.675 18.165 5.725 18.295 ;
		RECT	3.06 17.935 3.11 18.065 ;
		RECT	1.085 17.475 1.135 17.605 ;
		RECT	1.405 17.515 1.455 17.565 ;
		RECT	4.47 17.515 4.6 17.565 ;
		RECT	3.06 15.515 3.11 15.645 ;
		RECT	1.57 15.285 1.62 15.415 ;
		RECT	2.58 15.285 2.63 15.415 ;
		RECT	3.84 15.285 3.89 15.415 ;
		RECT	5.675 15.285 5.725 15.415 ;
		RECT	3.06 15.055 3.11 15.185 ;
		RECT	1.085 14.595 1.135 14.725 ;
		RECT	1.405 14.635 1.455 14.685 ;
		RECT	4.47 14.635 4.6 14.685 ;
		RECT	3.06 12.635 3.11 12.765 ;
		RECT	1.57 12.405 1.62 12.535 ;
		RECT	2.58 12.405 2.63 12.535 ;
		RECT	3.84 12.405 3.89 12.535 ;
		RECT	5.675 12.405 5.725 12.535 ;
		RECT	3.06 12.175 3.11 12.305 ;
		RECT	1.085 11.715 1.135 11.845 ;
		RECT	1.405 11.755 1.455 11.805 ;
		RECT	4.47 11.755 4.6 11.805 ;
		RECT	3.06 9.755 3.11 9.885 ;
		RECT	1.57 9.525 1.62 9.655 ;
		RECT	2.58 9.525 2.63 9.655 ;
		RECT	3.84 9.525 3.89 9.655 ;
		RECT	5.675 9.525 5.725 9.655 ;
		RECT	3.06 9.295 3.11 9.425 ;
		RECT	1.085 8.835 1.135 8.965 ;
		RECT	1.405 8.875 1.455 8.925 ;
		RECT	4.47 8.875 4.6 8.925 ;
		RECT	3.06 6.875 3.11 7.005 ;
		RECT	1.57 6.645 1.62 6.775 ;
		RECT	2.58 6.645 2.63 6.775 ;
		RECT	3.84 6.645 3.89 6.775 ;
		RECT	5.675 6.645 5.725 6.775 ;
		RECT	3.06 6.415 3.11 6.545 ;
		RECT	1.085 5.955 1.135 6.085 ;
		RECT	1.405 5.995 1.455 6.045 ;
		RECT	4.47 5.995 4.6 6.045 ;
		RECT	3.06 3.995 3.11 4.125 ;
		RECT	1.57 3.765 1.62 3.895 ;
		RECT	2.58 3.765 2.63 3.895 ;
		RECT	3.84 3.765 3.89 3.895 ;
		RECT	5.675 3.765 5.725 3.895 ;
		RECT	3.06 3.535 3.11 3.665 ;
		RECT	1.085 3.075 1.135 3.205 ;
		RECT	1.405 3.115 1.455 3.165 ;
		RECT	4.47 3.115 4.6 3.165 ;
		RECT	3.06 1.115 3.11 1.245 ;
		RECT	1.57 0.885 1.62 1.015 ;
		RECT	2.58 0.885 2.63 1.015 ;
		RECT	3.84 0.885 3.89 1.015 ;
		RECT	5.675 0.885 5.725 1.015 ;
		RECT	3.06 26.575 3.11 26.705 ;
		RECT	1.085 26.115 1.135 26.245 ;
		RECT	1.405 26.155 1.455 26.205 ;
		RECT	4.47 26.155 4.6 26.205 ;
		RECT	3.06 24.155 3.11 24.285 ;
		RECT	1.57 23.925 1.62 24.055 ;
		RECT	2.58 23.925 2.63 24.055 ;
		RECT	3.84 23.925 3.89 24.055 ;
		RECT	5.675 23.925 5.725 24.055 ;
		RECT	0.435 26.115 0.485 26.245 ;
		RECT	0.435 26.575 0.485 26.705 ;
		RECT	0.435 24.155 0.485 24.285 ;
		RECT	0.435 23.235 0.485 23.365 ;
		RECT	0.435 23.695 0.485 23.825 ;
		RECT	0.435 21.275 0.485 21.405 ;
		RECT	0.435 20.355 0.485 20.485 ;
		RECT	0.435 20.815 0.485 20.945 ;
		RECT	0.435 18.395 0.485 18.525 ;
		RECT	0.435 17.475 0.485 17.605 ;
		RECT	0.435 17.935 0.485 18.065 ;
		RECT	0.435 15.515 0.485 15.645 ;
		RECT	0.435 14.595 0.485 14.725 ;
		RECT	0.435 15.055 0.485 15.185 ;
		RECT	0.435 12.635 0.485 12.765 ;
		RECT	0.435 11.715 0.485 11.845 ;
		RECT	0.435 12.175 0.485 12.305 ;
		RECT	0.435 9.755 0.485 9.885 ;
		RECT	0.435 8.835 0.485 8.965 ;
		RECT	0.435 9.295 0.485 9.425 ;
		RECT	0.435 6.875 0.485 7.005 ;
		RECT	0.435 5.955 0.485 6.085 ;
		RECT	0.435 6.415 0.485 6.545 ;
		RECT	0.435 3.995 0.485 4.125 ;
		RECT	0.435 3.075 0.485 3.205 ;
		RECT	0.435 3.535 0.485 3.665 ;
		RECT	0.435 1.115 0.485 1.245 ;
		RECT	6.22 71.355 6.27 71.485 ;
		RECT	7.5 71.355 7.55 71.485 ;
		RECT	9.04 71.355 9.09 71.485 ;
		RECT	9.315 71.355 9.365 71.485 ;
		RECT	9.72 71.355 9.77 71.485 ;
		RECT	11.025 71.355 11.075 71.485 ;
		RECT	12.79 71.355 12.84 71.485 ;
		RECT	6.225 73.775 6.275 73.905 ;
		RECT	7.5 73.775 7.55 73.905 ;
		RECT	9.04 73.775 9.09 73.905 ;
		RECT	9.315 73.775 9.365 73.905 ;
		RECT	11.025 73.775 11.075 73.905 ;
		RECT	12.79 73.775 12.84 73.905 ;
		RECT	7.18 74.005 7.23 74.135 ;
		RECT	14.14 74.005 14.19 74.135 ;
		RECT	8.56 71.355 8.61 71.485 ;
		RECT	10.27 71.355 10.32 71.485 ;
		RECT	8.56 73.775 8.61 73.905 ;
		RECT	10.27 73.775 10.32 73.905 ;
		RECT	6.22 74.235 6.27 74.365 ;
		RECT	7.5 74.235 7.55 74.365 ;
		RECT	9.04 74.235 9.09 74.365 ;
		RECT	9.315 74.235 9.365 74.365 ;
		RECT	9.72 74.235 9.77 74.365 ;
		RECT	11.025 74.235 11.075 74.365 ;
		RECT	12.79 74.235 12.84 74.365 ;
		RECT	6.225 76.655 6.275 76.785 ;
		RECT	7.5 76.655 7.55 76.785 ;
		RECT	9.04 76.655 9.09 76.785 ;
		RECT	9.315 76.655 9.365 76.785 ;
		RECT	11.025 76.655 11.075 76.785 ;
		RECT	12.79 76.655 12.84 76.785 ;
		RECT	7.18 76.885 7.23 77.015 ;
		RECT	14.14 76.885 14.19 77.015 ;
		RECT	8.56 74.235 8.61 74.365 ;
		RECT	10.27 74.235 10.32 74.365 ;
		RECT	8.56 76.655 8.61 76.785 ;
		RECT	10.27 76.655 10.32 76.785 ;
		RECT	6.22 77.115 6.27 77.245 ;
		RECT	7.5 77.115 7.55 77.245 ;
		RECT	9.04 77.115 9.09 77.245 ;
		RECT	9.315 77.115 9.365 77.245 ;
		RECT	9.72 77.115 9.77 77.245 ;
		RECT	11.025 77.115 11.075 77.245 ;
		RECT	12.79 77.115 12.84 77.245 ;
		RECT	6.225 79.535 6.275 79.665 ;
		RECT	7.5 79.535 7.55 79.665 ;
		RECT	9.04 79.535 9.09 79.665 ;
		RECT	9.315 79.535 9.365 79.665 ;
		RECT	11.025 79.535 11.075 79.665 ;
		RECT	12.79 79.535 12.84 79.665 ;
		RECT	7.18 79.765 7.23 79.895 ;
		RECT	14.14 79.765 14.19 79.895 ;
		RECT	8.56 77.115 8.61 77.245 ;
		RECT	10.27 77.115 10.32 77.245 ;
		RECT	8.56 79.535 8.61 79.665 ;
		RECT	10.27 79.535 10.32 79.665 ;
		RECT	6.22 79.995 6.27 80.125 ;
		RECT	7.5 79.995 7.55 80.125 ;
		RECT	9.04 79.995 9.09 80.125 ;
		RECT	9.315 79.995 9.365 80.125 ;
		RECT	9.72 79.995 9.77 80.125 ;
		RECT	11.025 79.995 11.075 80.125 ;
		RECT	12.79 79.995 12.84 80.125 ;
		RECT	6.225 82.415 6.275 82.545 ;
		RECT	7.5 82.415 7.55 82.545 ;
		RECT	9.04 82.415 9.09 82.545 ;
		RECT	9.315 82.415 9.365 82.545 ;
		RECT	11.025 82.415 11.075 82.545 ;
		RECT	12.79 82.415 12.84 82.545 ;
		RECT	7.18 82.645 7.23 82.775 ;
		RECT	14.14 82.645 14.19 82.775 ;
		RECT	8.56 79.995 8.61 80.125 ;
		RECT	10.27 79.995 10.32 80.125 ;
		RECT	8.56 82.415 8.61 82.545 ;
		RECT	10.27 82.415 10.32 82.545 ;
		RECT	6.22 82.875 6.27 83.005 ;
		RECT	7.5 82.875 7.55 83.005 ;
		RECT	9.04 82.875 9.09 83.005 ;
		RECT	9.315 82.875 9.365 83.005 ;
		RECT	9.72 82.875 9.77 83.005 ;
		RECT	11.025 82.875 11.075 83.005 ;
		RECT	12.79 82.875 12.84 83.005 ;
		RECT	6.225 85.295 6.275 85.425 ;
		RECT	7.5 85.295 7.55 85.425 ;
		RECT	9.04 85.295 9.09 85.425 ;
		RECT	9.315 85.295 9.365 85.425 ;
		RECT	11.025 85.295 11.075 85.425 ;
		RECT	12.79 85.295 12.84 85.425 ;
		RECT	7.18 85.525 7.23 85.655 ;
		RECT	14.14 85.525 14.19 85.655 ;
		RECT	8.56 82.875 8.61 83.005 ;
		RECT	10.27 82.875 10.32 83.005 ;
		RECT	8.56 85.295 8.61 85.425 ;
		RECT	10.27 85.295 10.32 85.425 ;
		RECT	6.22 85.755 6.27 85.885 ;
		RECT	7.5 85.755 7.55 85.885 ;
		RECT	9.04 85.755 9.09 85.885 ;
		RECT	9.315 85.755 9.365 85.885 ;
		RECT	9.72 85.755 9.77 85.885 ;
		RECT	11.025 85.755 11.075 85.885 ;
		RECT	12.79 85.755 12.84 85.885 ;
		RECT	6.225 88.175 6.275 88.305 ;
		RECT	7.5 88.175 7.55 88.305 ;
		RECT	9.04 88.175 9.09 88.305 ;
		RECT	9.315 88.175 9.365 88.305 ;
		RECT	11.025 88.175 11.075 88.305 ;
		RECT	12.79 88.175 12.84 88.305 ;
		RECT	7.18 88.405 7.23 88.535 ;
		RECT	14.14 88.405 14.19 88.535 ;
		RECT	8.56 85.755 8.61 85.885 ;
		RECT	10.27 85.755 10.32 85.885 ;
		RECT	8.56 88.175 8.61 88.305 ;
		RECT	10.27 88.175 10.32 88.305 ;
		RECT	6.22 88.635 6.27 88.765 ;
		RECT	7.5 88.635 7.55 88.765 ;
		RECT	9.04 88.635 9.09 88.765 ;
		RECT	9.315 88.635 9.365 88.765 ;
		RECT	9.72 88.635 9.77 88.765 ;
		RECT	11.025 88.635 11.075 88.765 ;
		RECT	12.79 88.635 12.84 88.765 ;
		RECT	6.225 91.055 6.275 91.185 ;
		RECT	7.5 91.055 7.55 91.185 ;
		RECT	9.04 91.055 9.09 91.185 ;
		RECT	9.315 91.055 9.365 91.185 ;
		RECT	11.025 91.055 11.075 91.185 ;
		RECT	12.79 91.055 12.84 91.185 ;
		RECT	7.18 91.285 7.23 91.415 ;
		RECT	14.14 91.285 14.19 91.415 ;
		RECT	8.56 88.635 8.61 88.765 ;
		RECT	10.27 88.635 10.32 88.765 ;
		RECT	8.56 91.055 8.61 91.185 ;
		RECT	10.27 91.055 10.32 91.185 ;
		RECT	6.22 91.515 6.27 91.645 ;
		RECT	7.5 91.515 7.55 91.645 ;
		RECT	9.04 91.515 9.09 91.645 ;
		RECT	9.315 91.515 9.365 91.645 ;
		RECT	9.72 91.515 9.77 91.645 ;
		RECT	11.025 91.515 11.075 91.645 ;
		RECT	12.79 91.515 12.84 91.645 ;
		RECT	6.225 93.935 6.275 94.065 ;
		RECT	7.5 93.935 7.55 94.065 ;
		RECT	9.04 93.935 9.09 94.065 ;
		RECT	9.315 93.935 9.365 94.065 ;
		RECT	11.025 93.935 11.075 94.065 ;
		RECT	12.79 93.935 12.84 94.065 ;
		RECT	7.18 94.165 7.23 94.295 ;
		RECT	14.14 94.165 14.19 94.295 ;
		RECT	8.56 91.515 8.61 91.645 ;
		RECT	10.27 91.515 10.32 91.645 ;
		RECT	8.56 93.935 8.61 94.065 ;
		RECT	10.27 93.935 10.32 94.065 ;
		RECT	6.22 94.395 6.27 94.525 ;
		RECT	7.5 94.395 7.55 94.525 ;
		RECT	9.04 94.395 9.09 94.525 ;
		RECT	9.315 94.395 9.365 94.525 ;
		RECT	9.72 94.395 9.77 94.525 ;
		RECT	11.025 94.395 11.075 94.525 ;
		RECT	12.79 94.395 12.84 94.525 ;
		RECT	6.225 96.815 6.275 96.945 ;
		RECT	7.5 96.815 7.55 96.945 ;
		RECT	9.04 96.815 9.09 96.945 ;
		RECT	9.315 96.815 9.365 96.945 ;
		RECT	11.025 96.815 11.075 96.945 ;
		RECT	12.79 96.815 12.84 96.945 ;
		RECT	7.18 97.045 7.23 97.175 ;
		RECT	14.14 97.045 14.19 97.175 ;
		RECT	8.56 94.395 8.61 94.525 ;
		RECT	10.27 94.395 10.32 94.525 ;
		RECT	8.56 96.815 8.61 96.945 ;
		RECT	10.27 96.815 10.32 96.945 ;
		RECT	6.22 97.275 6.27 97.405 ;
		RECT	7.5 97.275 7.55 97.405 ;
		RECT	9.04 97.275 9.09 97.405 ;
		RECT	9.315 97.275 9.365 97.405 ;
		RECT	9.72 97.275 9.77 97.405 ;
		RECT	11.025 97.275 11.075 97.405 ;
		RECT	12.79 97.275 12.84 97.405 ;
		RECT	6.225 99.695 6.275 99.825 ;
		RECT	7.5 99.695 7.55 99.825 ;
		RECT	9.04 99.695 9.09 99.825 ;
		RECT	9.315 99.695 9.365 99.825 ;
		RECT	11.025 99.695 11.075 99.825 ;
		RECT	12.79 99.695 12.84 99.825 ;
		RECT	7.18 99.925 7.23 100.055 ;
		RECT	14.14 99.925 14.19 100.055 ;
		RECT	8.56 97.275 8.61 97.405 ;
		RECT	10.27 97.275 10.32 97.405 ;
		RECT	8.56 99.695 8.61 99.825 ;
		RECT	10.27 99.695 10.32 99.825 ;
		RECT	14.33 74.235 14.38 74.365 ;
		RECT	6.22 74.695 6.27 74.825 ;
		RECT	7.5 74.695 7.55 74.825 ;
		RECT	9.04 74.695 9.09 74.825 ;
		RECT	9.315 74.695 9.365 74.825 ;
		RECT	9.72 74.695 9.77 74.825 ;
		RECT	11.025 74.695 11.075 74.825 ;
		RECT	12.79 74.695 12.84 74.825 ;
		RECT	14.33 76.655 14.38 76.785 ;
		RECT	5.675 76.885 5.725 77.015 ;
		RECT	6.065 76.885 6.115 77.015 ;
		RECT	6.725 76.885 6.775 77.015 ;
		RECT	8.42 76.885 8.47 77.015 ;
		RECT	8.77 76.885 8.82 77.015 ;
		RECT	11.555 76.885 11.605 77.015 ;
		RECT	11.815 76.885 11.865 77.015 ;
		RECT	12.52 76.885 12.57 77.015 ;
		RECT	13.98 76.885 14.03 77.015 ;
		RECT	14.33 77.115 14.38 77.245 ;
		RECT	6.22 77.575 6.27 77.705 ;
		RECT	7.5 77.575 7.55 77.705 ;
		RECT	9.04 77.575 9.09 77.705 ;
		RECT	9.315 77.575 9.365 77.705 ;
		RECT	9.72 77.575 9.77 77.705 ;
		RECT	11.025 77.575 11.075 77.705 ;
		RECT	12.79 77.575 12.84 77.705 ;
		RECT	14.33 79.535 14.38 79.665 ;
		RECT	5.675 79.765 5.725 79.895 ;
		RECT	6.065 79.765 6.115 79.895 ;
		RECT	6.725 79.765 6.775 79.895 ;
		RECT	8.42 79.765 8.47 79.895 ;
		RECT	8.77 79.765 8.82 79.895 ;
		RECT	11.555 79.765 11.605 79.895 ;
		RECT	11.815 79.765 11.865 79.895 ;
		RECT	12.52 79.765 12.57 79.895 ;
		RECT	13.98 79.765 14.03 79.895 ;
		RECT	14.33 79.995 14.38 80.125 ;
		RECT	6.22 80.455 6.27 80.585 ;
		RECT	7.5 80.455 7.55 80.585 ;
		RECT	9.04 80.455 9.09 80.585 ;
		RECT	9.315 80.455 9.365 80.585 ;
		RECT	9.72 80.455 9.77 80.585 ;
		RECT	11.025 80.455 11.075 80.585 ;
		RECT	12.79 80.455 12.84 80.585 ;
		RECT	14.33 82.415 14.38 82.545 ;
		RECT	5.675 82.645 5.725 82.775 ;
		RECT	6.065 82.645 6.115 82.775 ;
		RECT	6.725 82.645 6.775 82.775 ;
		RECT	8.42 82.645 8.47 82.775 ;
		RECT	8.77 82.645 8.82 82.775 ;
		RECT	11.555 82.645 11.605 82.775 ;
		RECT	11.815 82.645 11.865 82.775 ;
		RECT	12.52 82.645 12.57 82.775 ;
		RECT	13.98 82.645 14.03 82.775 ;
		RECT	14.33 82.875 14.38 83.005 ;
		RECT	6.22 83.335 6.27 83.465 ;
		RECT	7.5 83.335 7.55 83.465 ;
		RECT	9.04 83.335 9.09 83.465 ;
		RECT	9.315 83.335 9.365 83.465 ;
		RECT	9.72 83.335 9.77 83.465 ;
		RECT	11.025 83.335 11.075 83.465 ;
		RECT	12.79 83.335 12.84 83.465 ;
		RECT	14.33 85.295 14.38 85.425 ;
		RECT	5.675 85.525 5.725 85.655 ;
		RECT	6.065 85.525 6.115 85.655 ;
		RECT	6.725 85.525 6.775 85.655 ;
		RECT	8.42 85.525 8.47 85.655 ;
		RECT	8.77 85.525 8.82 85.655 ;
		RECT	11.555 85.525 11.605 85.655 ;
		RECT	11.815 85.525 11.865 85.655 ;
		RECT	12.52 85.525 12.57 85.655 ;
		RECT	13.98 85.525 14.03 85.655 ;
		RECT	14.33 85.755 14.38 85.885 ;
		RECT	6.22 86.215 6.27 86.345 ;
		RECT	7.5 86.215 7.55 86.345 ;
		RECT	9.04 86.215 9.09 86.345 ;
		RECT	9.315 86.215 9.365 86.345 ;
		RECT	9.72 86.215 9.77 86.345 ;
		RECT	11.025 86.215 11.075 86.345 ;
		RECT	12.79 86.215 12.84 86.345 ;
		RECT	14.33 88.175 14.38 88.305 ;
		RECT	5.675 88.405 5.725 88.535 ;
		RECT	6.065 88.405 6.115 88.535 ;
		RECT	6.725 88.405 6.775 88.535 ;
		RECT	8.42 88.405 8.47 88.535 ;
		RECT	8.77 88.405 8.82 88.535 ;
		RECT	11.555 88.405 11.605 88.535 ;
		RECT	11.815 88.405 11.865 88.535 ;
		RECT	12.52 88.405 12.57 88.535 ;
		RECT	13.98 88.405 14.03 88.535 ;
		RECT	14.33 88.635 14.38 88.765 ;
		RECT	6.22 89.095 6.27 89.225 ;
		RECT	7.5 89.095 7.55 89.225 ;
		RECT	9.04 89.095 9.09 89.225 ;
		RECT	9.315 89.095 9.365 89.225 ;
		RECT	9.72 89.095 9.77 89.225 ;
		RECT	11.025 89.095 11.075 89.225 ;
		RECT	12.79 89.095 12.84 89.225 ;
		RECT	14.33 91.055 14.38 91.185 ;
		RECT	5.675 91.285 5.725 91.415 ;
		RECT	6.065 91.285 6.115 91.415 ;
		RECT	6.725 91.285 6.775 91.415 ;
		RECT	8.42 91.285 8.47 91.415 ;
		RECT	8.77 91.285 8.82 91.415 ;
		RECT	11.555 91.285 11.605 91.415 ;
		RECT	11.815 91.285 11.865 91.415 ;
		RECT	12.52 91.285 12.57 91.415 ;
		RECT	13.98 91.285 14.03 91.415 ;
		RECT	14.33 91.515 14.38 91.645 ;
		RECT	6.22 91.975 6.27 92.105 ;
		RECT	7.5 91.975 7.55 92.105 ;
		RECT	9.04 91.975 9.09 92.105 ;
		RECT	9.315 91.975 9.365 92.105 ;
		RECT	9.72 91.975 9.77 92.105 ;
		RECT	11.025 91.975 11.075 92.105 ;
		RECT	12.79 91.975 12.84 92.105 ;
		RECT	14.33 93.935 14.38 94.065 ;
		RECT	5.675 94.165 5.725 94.295 ;
		RECT	6.065 94.165 6.115 94.295 ;
		RECT	6.725 94.165 6.775 94.295 ;
		RECT	8.42 94.165 8.47 94.295 ;
		RECT	8.77 94.165 8.82 94.295 ;
		RECT	11.555 94.165 11.605 94.295 ;
		RECT	11.815 94.165 11.865 94.295 ;
		RECT	12.52 94.165 12.57 94.295 ;
		RECT	13.98 94.165 14.03 94.295 ;
		RECT	14.33 94.395 14.38 94.525 ;
		RECT	6.22 94.855 6.27 94.985 ;
		RECT	7.5 94.855 7.55 94.985 ;
		RECT	9.04 94.855 9.09 94.985 ;
		RECT	9.315 94.855 9.365 94.985 ;
		RECT	9.72 94.855 9.77 94.985 ;
		RECT	11.025 94.855 11.075 94.985 ;
		RECT	12.79 94.855 12.84 94.985 ;
		RECT	14.33 96.815 14.38 96.945 ;
		RECT	5.675 97.045 5.725 97.175 ;
		RECT	6.065 97.045 6.115 97.175 ;
		RECT	6.725 97.045 6.775 97.175 ;
		RECT	8.42 97.045 8.47 97.175 ;
		RECT	8.77 97.045 8.82 97.175 ;
		RECT	11.555 97.045 11.605 97.175 ;
		RECT	11.815 97.045 11.865 97.175 ;
		RECT	12.52 97.045 12.57 97.175 ;
		RECT	13.98 97.045 14.03 97.175 ;
		RECT	14.33 97.275 14.38 97.405 ;
		RECT	6.22 97.735 6.27 97.865 ;
		RECT	7.5 97.735 7.55 97.865 ;
		RECT	9.04 97.735 9.09 97.865 ;
		RECT	9.315 97.735 9.365 97.865 ;
		RECT	9.72 97.735 9.77 97.865 ;
		RECT	11.025 97.735 11.075 97.865 ;
		RECT	12.79 97.735 12.84 97.865 ;
		RECT	14.33 99.695 14.38 99.825 ;
		RECT	5.675 99.925 5.725 100.055 ;
		RECT	6.065 99.925 6.115 100.055 ;
		RECT	6.725 99.925 6.775 100.055 ;
		RECT	8.42 99.925 8.47 100.055 ;
		RECT	8.77 99.925 8.82 100.055 ;
		RECT	11.555 99.925 11.605 100.055 ;
		RECT	11.815 99.925 11.865 100.055 ;
		RECT	12.52 99.925 12.57 100.055 ;
		RECT	13.98 99.925 14.03 100.055 ;
		RECT	14.33 71.355 14.38 71.485 ;
		RECT	6.22 71.815 6.27 71.945 ;
		RECT	7.5 71.815 7.55 71.945 ;
		RECT	9.04 71.815 9.09 71.945 ;
		RECT	9.315 71.815 9.365 71.945 ;
		RECT	9.72 71.815 9.77 71.945 ;
		RECT	11.025 71.815 11.075 71.945 ;
		RECT	12.79 71.815 12.84 71.945 ;
		RECT	14.33 73.775 14.38 73.905 ;
		RECT	5.675 74.005 5.725 74.135 ;
		RECT	6.065 74.005 6.115 74.135 ;
		RECT	6.725 74.005 6.775 74.135 ;
		RECT	8.42 74.005 8.47 74.135 ;
		RECT	8.77 74.005 8.82 74.135 ;
		RECT	11.555 74.005 11.605 74.135 ;
		RECT	11.815 74.005 11.865 74.135 ;
		RECT	12.52 74.005 12.57 74.135 ;
		RECT	13.98 74.005 14.03 74.135 ;
		RECT	13.98 100.615 14.03 100.745 ;
		RECT	1.57 100.615 1.62 100.745 ;
		RECT	2.485 100.615 2.665 100.745 ;
		RECT	3.84 100.615 3.89 100.745 ;
		RECT	7.19 100.615 7.24 100.745 ;
		RECT	14.14 100.615 14.19 100.745 ;
		RECT	13.8 100.385 13.85 100.515 ;
		RECT	8.56 100.155 8.61 100.285 ;
		RECT	10.27 100.155 10.32 100.285 ;
		RECT	0.435 100.155 0.485 100.285 ;
		RECT	0.62 100.615 0.67 100.745 ;
		RECT	3.65 100.615 3.7 100.745 ;
		RECT	2.18 100.155 2.23 100.285 ;
		RECT	0.9 76.885 0.95 77.015 ;
		RECT	0.9 79.765 0.95 79.895 ;
		RECT	0.9 82.645 0.95 82.775 ;
		RECT	0.9 85.525 0.95 85.655 ;
		RECT	0.9 88.405 0.95 88.535 ;
		RECT	0.9 91.285 0.95 91.415 ;
		RECT	0.9 94.165 0.95 94.295 ;
		RECT	0.9 97.045 0.95 97.175 ;
		RECT	0.9 99.925 0.95 100.055 ;
		RECT	0.9 74.005 0.95 74.135 ;
		RECT	3.65 74.005 3.7 74.135 ;
		RECT	3.65 76.885 3.7 77.015 ;
		RECT	3.65 79.765 3.7 79.895 ;
		RECT	3.65 82.645 3.7 82.775 ;
		RECT	3.65 85.525 3.7 85.655 ;
		RECT	3.65 88.405 3.7 88.535 ;
		RECT	3.65 91.285 3.7 91.415 ;
		RECT	3.65 94.165 3.7 94.295 ;
		RECT	3.65 97.045 3.7 97.175 ;
		RECT	3.65 99.925 3.7 100.055 ;
		RECT	2.18 71.355 2.23 71.485 ;
		RECT	2.18 73.775 2.23 73.905 ;
		RECT	2.18 74.235 2.23 74.365 ;
		RECT	2.18 76.655 2.23 76.785 ;
		RECT	2.18 77.115 2.23 77.245 ;
		RECT	2.18 79.535 2.23 79.665 ;
		RECT	2.18 79.995 2.23 80.125 ;
		RECT	2.18 82.415 2.23 82.545 ;
		RECT	2.18 82.875 2.23 83.005 ;
		RECT	2.18 85.295 2.23 85.425 ;
		RECT	2.18 85.755 2.23 85.885 ;
		RECT	2.18 88.175 2.23 88.305 ;
		RECT	2.18 88.635 2.23 88.765 ;
		RECT	2.18 91.055 2.23 91.185 ;
		RECT	2.18 91.515 2.23 91.645 ;
		RECT	2.18 93.935 2.23 94.065 ;
		RECT	2.18 94.395 2.23 94.525 ;
		RECT	2.18 96.815 2.23 96.945 ;
		RECT	2.18 97.275 2.23 97.405 ;
		RECT	2.18 99.695 2.23 99.825 ;
		RECT	3.06 74.235 3.11 74.365 ;
		RECT	1.085 74.695 1.135 74.825 ;
		RECT	1.405 74.735 1.455 74.785 ;
		RECT	4.47 74.735 4.6 74.785 ;
		RECT	3.06 76.655 3.11 76.785 ;
		RECT	1.57 76.885 1.62 77.015 ;
		RECT	2.58 76.885 2.63 77.015 ;
		RECT	3.84 76.885 3.89 77.015 ;
		RECT	5.675 76.885 5.725 77.015 ;
		RECT	3.06 77.115 3.11 77.245 ;
		RECT	1.085 77.575 1.135 77.705 ;
		RECT	1.405 77.615 1.455 77.665 ;
		RECT	4.47 77.615 4.6 77.665 ;
		RECT	3.06 79.535 3.11 79.665 ;
		RECT	1.57 79.765 1.62 79.895 ;
		RECT	2.58 79.765 2.63 79.895 ;
		RECT	3.84 79.765 3.89 79.895 ;
		RECT	5.675 79.765 5.725 79.895 ;
		RECT	3.06 79.995 3.11 80.125 ;
		RECT	1.085 80.455 1.135 80.585 ;
		RECT	1.405 80.495 1.455 80.545 ;
		RECT	4.47 80.495 4.6 80.545 ;
		RECT	3.06 82.415 3.11 82.545 ;
		RECT	1.57 82.645 1.62 82.775 ;
		RECT	2.58 82.645 2.63 82.775 ;
		RECT	3.84 82.645 3.89 82.775 ;
		RECT	5.675 82.645 5.725 82.775 ;
		RECT	3.06 82.875 3.11 83.005 ;
		RECT	1.085 83.335 1.135 83.465 ;
		RECT	1.405 83.375 1.455 83.425 ;
		RECT	4.47 83.375 4.6 83.425 ;
		RECT	3.06 85.295 3.11 85.425 ;
		RECT	1.57 85.525 1.62 85.655 ;
		RECT	2.58 85.525 2.63 85.655 ;
		RECT	3.84 85.525 3.89 85.655 ;
		RECT	5.675 85.525 5.725 85.655 ;
		RECT	3.06 85.755 3.11 85.885 ;
		RECT	1.085 86.215 1.135 86.345 ;
		RECT	1.405 86.255 1.455 86.305 ;
		RECT	4.47 86.255 4.6 86.305 ;
		RECT	3.06 88.175 3.11 88.305 ;
		RECT	1.57 88.405 1.62 88.535 ;
		RECT	2.58 88.405 2.63 88.535 ;
		RECT	3.84 88.405 3.89 88.535 ;
		RECT	5.675 88.405 5.725 88.535 ;
		RECT	3.06 88.635 3.11 88.765 ;
		RECT	1.085 89.095 1.135 89.225 ;
		RECT	1.405 89.135 1.455 89.185 ;
		RECT	4.47 89.135 4.6 89.185 ;
		RECT	3.06 91.055 3.11 91.185 ;
		RECT	1.57 91.285 1.62 91.415 ;
		RECT	2.58 91.285 2.63 91.415 ;
		RECT	3.84 91.285 3.89 91.415 ;
		RECT	5.675 91.285 5.725 91.415 ;
		RECT	3.06 91.515 3.11 91.645 ;
		RECT	1.085 91.975 1.135 92.105 ;
		RECT	1.405 92.015 1.455 92.065 ;
		RECT	4.47 92.015 4.6 92.065 ;
		RECT	3.06 93.935 3.11 94.065 ;
		RECT	1.57 94.165 1.62 94.295 ;
		RECT	2.58 94.165 2.63 94.295 ;
		RECT	3.84 94.165 3.89 94.295 ;
		RECT	5.675 94.165 5.725 94.295 ;
		RECT	3.06 94.395 3.11 94.525 ;
		RECT	1.085 94.855 1.135 94.985 ;
		RECT	1.405 94.895 1.455 94.945 ;
		RECT	4.47 94.895 4.6 94.945 ;
		RECT	3.06 96.815 3.11 96.945 ;
		RECT	1.57 97.045 1.62 97.175 ;
		RECT	2.58 97.045 2.63 97.175 ;
		RECT	3.84 97.045 3.89 97.175 ;
		RECT	5.675 97.045 5.725 97.175 ;
		RECT	3.06 97.275 3.11 97.405 ;
		RECT	1.085 97.735 1.135 97.865 ;
		RECT	1.405 97.775 1.455 97.825 ;
		RECT	4.47 97.775 4.6 97.825 ;
		RECT	3.06 99.695 3.11 99.825 ;
		RECT	1.57 99.925 1.62 100.055 ;
		RECT	2.58 99.925 2.63 100.055 ;
		RECT	3.84 99.925 3.89 100.055 ;
		RECT	5.675 99.925 5.725 100.055 ;
		RECT	3.06 71.355 3.11 71.485 ;
		RECT	1.085 71.815 1.135 71.945 ;
		RECT	1.405 71.855 1.455 71.905 ;
		RECT	4.47 71.855 4.6 71.905 ;
		RECT	3.06 73.775 3.11 73.905 ;
		RECT	1.57 74.005 1.62 74.135 ;
		RECT	2.58 74.005 2.63 74.135 ;
		RECT	3.84 74.005 3.89 74.135 ;
		RECT	5.675 74.005 5.725 74.135 ;
		RECT	0.435 71.815 0.485 71.945 ;
		RECT	0.435 71.355 0.485 71.485 ;
		RECT	0.435 73.775 0.485 73.905 ;
		RECT	0.435 74.695 0.485 74.825 ;
		RECT	0.435 74.235 0.485 74.365 ;
		RECT	0.435 76.655 0.485 76.785 ;
		RECT	0.435 77.575 0.485 77.705 ;
		RECT	0.435 77.115 0.485 77.245 ;
		RECT	0.435 79.535 0.485 79.665 ;
		RECT	0.435 80.455 0.485 80.585 ;
		RECT	0.435 79.995 0.485 80.125 ;
		RECT	0.435 82.415 0.485 82.545 ;
		RECT	0.435 83.335 0.485 83.465 ;
		RECT	0.435 82.875 0.485 83.005 ;
		RECT	0.435 85.295 0.485 85.425 ;
		RECT	0.435 86.215 0.485 86.345 ;
		RECT	0.435 85.755 0.485 85.885 ;
		RECT	0.435 88.175 0.485 88.305 ;
		RECT	0.435 89.095 0.485 89.225 ;
		RECT	0.435 88.635 0.485 88.765 ;
		RECT	0.435 91.055 0.485 91.185 ;
		RECT	0.435 91.975 0.485 92.105 ;
		RECT	0.435 91.515 0.485 91.645 ;
		RECT	0.435 93.935 0.485 94.065 ;
		RECT	0.435 94.855 0.485 94.985 ;
		RECT	0.435 94.395 0.485 94.525 ;
		RECT	0.435 96.815 0.485 96.945 ;
		RECT	0.435 97.735 0.485 97.865 ;
		RECT	0.435 97.275 0.485 97.405 ;
		RECT	0.435 99.695 0.485 99.825 ;
		RECT	50.325 28.475 50.505 28.605 ;
		RECT	50.32 34.46 50.45 34.64 ;
		RECT	50.32 63.49 50.45 63.67 ;
		RECT	50.325 69.455 50.505 69.585 ;
		RECT	50.635 30.055 50.815 30.185 ;
		RECT	50.77 32.06 50.82 32.19 ;
		RECT	50.77 34.975 50.82 35.105 ;
		RECT	50.77 35.96 50.82 36.09 ;
		RECT	50.77 37.93 50.82 38.06 ;
		RECT	50.77 38.91 50.82 39.04 ;
		RECT	50.77 39.895 50.82 40.025 ;
		RECT	50.77 42.85 50.82 42.98 ;
		RECT	50.77 50.23 50.82 50.36 ;
		RECT	50.77 51.21 50.82 51.34 ;
		RECT	50.77 55.15 50.82 55.28 ;
		RECT	50.77 58.1 50.82 58.23 ;
		RECT	50.77 59.085 50.82 59.215 ;
		RECT	50.77 60.07 50.82 60.2 ;
		RECT	50.77 62.035 50.82 62.165 ;
		RECT	50.77 63.02 50.82 63.15 ;
		RECT	50.77 65.94 50.82 66.07 ;
		RECT	50.635 67.94 50.815 68.07 ;
		RECT	51.115 28.705 51.295 28.835 ;
		RECT	51.115 69.225 51.295 69.355 ;
		RECT	50.325 29.18 50.505 29.31 ;
		RECT	50.35 68.72 50.48 68.9 ;
		RECT	50.36 31.515 50.41 31.645 ;
		RECT	50.36 35.47 50.41 35.6 ;
		RECT	50.36 39.405 50.41 39.535 ;
		RECT	50.36 43.34 50.41 43.47 ;
		RECT	50.36 47.275 50.41 47.405 ;
		RECT	50.36 50.72 50.41 50.85 ;
		RECT	50.36 54.655 50.41 54.785 ;
		RECT	50.36 58.595 50.41 58.725 ;
		RECT	50.36 62.53 50.41 62.66 ;
		RECT	50.36 66.48 50.41 66.61 ;
		RECT	14.965 28.475 15.015 28.605 ;
		RECT	49.725 28.475 49.775 28.605 ;
		RECT	14.765 28.475 14.815 28.605 ;
		RECT	49.925 28.475 49.975 28.605 ;
		RECT	14.965 69.455 15.015 69.585 ;
		RECT	49.725 69.455 49.775 69.585 ;
		RECT	14.765 69.455 14.815 69.585 ;
		RECT	49.925 69.455 49.975 69.585 ;
		RECT	50.635 28.245 50.815 28.375 ;
		RECT	50.94 28.705 50.99 28.835 ;
		RECT	50.325 29.565 50.505 29.695 ;
		RECT	51.14 30.34 51.27 30.39 ;
		RECT	50.325 30.545 50.505 30.675 ;
		RECT	50.63 31.04 50.68 31.17 ;
		RECT	51.14 31.32 51.27 31.37 ;
		RECT	50.925 31.79 50.975 31.92 ;
		RECT	50.575 31.79 50.625 31.92 ;
		RECT	50.36 32.515 50.41 32.645 ;
		RECT	51.115 33.01 51.295 33.14 ;
		RECT	50.36 33.5 50.41 33.63 ;
		RECT	50.32 33.785 50.45 33.835 ;
		RECT	51.115 33.99 51.295 34.12 ;
		RECT	50.36 36.455 50.41 36.585 ;
		RECT	51.115 36.945 51.295 37.075 ;
		RECT	50.36 37.435 50.41 37.565 ;
		RECT	50.36 38.42 50.41 38.55 ;
		RECT	50.36 40.39 50.41 40.52 ;
		RECT	51.115 40.88 51.295 41.01 ;
		RECT	50.36 41.37 50.41 41.5 ;
		RECT	51.115 41.865 51.295 41.995 ;
		RECT	50.36 42.355 50.41 42.485 ;
		RECT	50.77 43.835 50.82 43.965 ;
		RECT	50.36 44.33 50.41 44.46 ;
		RECT	51.115 44.815 51.295 44.945 ;
		RECT	50.36 45.31 50.41 45.44 ;
		RECT	50.745 45.785 50.795 45.915 ;
		RECT	50.925 46.095 50.975 46.225 ;
		RECT	50.575 46.095 50.625 46.225 ;
		RECT	50.585 46.41 50.635 46.54 ;
		RECT	51.14 47.07 51.27 47.12 ;
		RECT	51.14 47.565 51.27 47.615 ;
		RECT	50.36 48.26 50.41 48.39 ;
		RECT	51.115 48.75 51.295 48.88 ;
		RECT	51.115 49.245 51.295 49.375 ;
		RECT	50.36 49.735 50.41 49.865 ;
		RECT	51.14 50.515 51.27 50.565 ;
		RECT	51.14 51.005 51.27 51.055 ;
		RECT	50.585 51.525 50.635 51.655 ;
		RECT	50.925 51.87 50.975 52 ;
		RECT	50.575 51.87 50.625 52 ;
		RECT	50.36 52.685 50.41 52.815 ;
		RECT	51.115 53.18 51.295 53.31 ;
		RECT	50.36 53.675 50.41 53.805 ;
		RECT	50.77 54.165 50.82 54.295 ;
		RECT	50.36 55.64 50.41 55.77 ;
		RECT	51.115 56.135 51.295 56.265 ;
		RECT	50.36 56.625 50.41 56.755 ;
		RECT	51.115 57.115 51.295 57.245 ;
		RECT	50.36 57.61 50.41 57.74 ;
		RECT	50.36 59.575 50.41 59.705 ;
		RECT	50.36 60.56 50.41 60.69 ;
		RECT	51.115 61.055 51.295 61.185 ;
		RECT	50.36 61.545 50.41 61.675 ;
		RECT	50.32 62.32 50.45 62.37 ;
		RECT	50.32 63.8 50.45 63.85 ;
		RECT	51.115 64.005 51.295 64.135 ;
		RECT	50.32 64.29 50.45 64.34 ;
		RECT	50.36 64.495 50.41 64.625 ;
		RECT	51.115 64.955 51.295 65.085 ;
		RECT	50.36 65.48 50.41 65.61 ;
		RECT	50.925 66.21 50.975 66.34 ;
		RECT	50.575 66.21 50.625 66.34 ;
		RECT	51.14 66.755 51.27 66.805 ;
		RECT	50.63 66.955 50.68 67.085 ;
		RECT	50.325 67.45 50.505 67.58 ;
		RECT	51.14 67.735 51.27 67.785 ;
		RECT	50.325 68.435 50.505 68.565 ;
		RECT	50.94 69.225 50.99 69.355 ;
		RECT	50.635 69.685 50.815 69.815 ;
		RECT	14.965 29.18 15.015 29.31 ;
		RECT	14.99 32.515 15.04 32.645 ;
		RECT	14.99 33.5 15.04 33.63 ;
		RECT	14.99 33.785 15.04 33.835 ;
		RECT	14.74 35.47 14.79 35.6 ;
		RECT	14.99 36.455 15.04 36.585 ;
		RECT	14.99 37.435 15.04 37.565 ;
		RECT	14.99 38.42 15.04 38.55 ;
		RECT	14.99 40.39 15.04 40.52 ;
		RECT	14.99 41.37 15.04 41.5 ;
		RECT	14.99 42.355 15.04 42.485 ;
		RECT	14.99 44.33 15.04 44.46 ;
		RECT	14.99 45.31 15.04 45.44 ;
		RECT	14.965 48.26 15.015 48.39 ;
		RECT	14.965 49.735 15.015 49.865 ;
		RECT	14.99 52.685 15.04 52.815 ;
		RECT	14.99 53.675 15.04 53.805 ;
		RECT	14.735 54.655 14.785 54.785 ;
		RECT	14.99 55.64 15.04 55.77 ;
		RECT	14.99 56.625 15.04 56.755 ;
		RECT	14.99 57.61 15.04 57.74 ;
		RECT	14.99 59.575 15.04 59.705 ;
		RECT	14.99 60.56 15.04 60.69 ;
		RECT	14.99 61.545 15.04 61.675 ;
		RECT	14.99 62.32 15.04 62.37 ;
		RECT	14.74 62.53 14.79 62.66 ;
		RECT	14.99 64.495 15.04 64.625 ;
		RECT	14.99 65.48 15.04 65.61 ;
		RECT	14.965 68.745 15.015 68.875 ;
		RECT	49.725 29.18 49.775 29.31 ;
		RECT	49.705 43.315 49.835 43.495 ;
		RECT	49.705 54.63 49.835 54.81 ;
		RECT	49.705 62.505 49.835 62.685 ;
		RECT	49.725 68.745 49.775 68.875 ;
		RECT	50.115 45.785 50.165 45.915 ;
		RECT	50.115 52.21 50.165 52.34 ;
		RECT	49.94 29.565 49.99 29.695 ;
		RECT	49.94 30.545 49.99 30.675 ;
		RECT	49.94 32.515 49.99 32.645 ;
		RECT	49.94 33.5 49.99 33.63 ;
		RECT	49.94 33.785 49.99 33.835 ;
		RECT	49.94 36.455 49.99 36.585 ;
		RECT	49.94 37.435 49.99 37.565 ;
		RECT	49.94 38.42 49.99 38.55 ;
		RECT	49.94 40.39 49.99 40.52 ;
		RECT	49.94 41.37 49.99 41.5 ;
		RECT	49.94 42.355 49.99 42.485 ;
		RECT	49.94 44.33 49.99 44.46 ;
		RECT	49.94 45.31 49.99 45.44 ;
		RECT	49.94 48.26 49.99 48.39 ;
		RECT	49.94 49.735 49.99 49.865 ;
		RECT	49.94 52.685 49.99 52.815 ;
		RECT	49.94 53.675 49.99 53.805 ;
		RECT	49.94 55.64 49.99 55.77 ;
		RECT	49.94 56.625 49.99 56.755 ;
		RECT	49.94 57.61 49.99 57.74 ;
		RECT	49.94 59.575 49.99 59.705 ;
		RECT	49.94 60.56 49.99 60.69 ;
		RECT	49.94 61.545 49.99 61.675 ;
		RECT	49.94 62.32 49.99 62.37 ;
		RECT	49.705 63.49 49.835 63.67 ;
		RECT	49.94 64.495 49.99 64.625 ;
		RECT	49.94 65.48 49.99 65.61 ;
		RECT	49.94 67.45 49.99 67.58 ;
		RECT	49.94 68.435 49.99 68.565 ;
		RECT	14.765 29.565 14.815 29.695 ;
		RECT	14.765 30.545 14.815 30.675 ;
		RECT	14.74 32.515 14.79 32.645 ;
		RECT	14.74 33.5 14.79 33.63 ;
		RECT	14.74 33.785 14.79 33.835 ;
		RECT	14.74 37.435 14.79 37.565 ;
		RECT	14.74 38.42 14.79 38.55 ;
		RECT	14.74 40.39 14.79 40.52 ;
		RECT	14.73 44.33 14.78 44.46 ;
		RECT	14.73 45.31 14.78 45.44 ;
		RECT	14.75 48.26 14.8 48.39 ;
		RECT	14.75 49.735 14.8 49.865 ;
		RECT	14.735 52.685 14.785 52.815 ;
		RECT	14.74 57.61 14.79 57.74 ;
		RECT	14.74 59.575 14.79 59.705 ;
		RECT	14.74 60.56 14.79 60.69 ;
		RECT	14.74 64.495 14.79 64.625 ;
		RECT	14.74 65.48 14.79 65.61 ;
		RECT	14.765 67.45 14.815 67.58 ;
		RECT	14.765 68.435 14.815 68.565 ;
		RECT	14.565 45.785 14.615 45.915 ;
		RECT	14.565 52.21 14.615 52.34 ;
		RECT	23.975 43.835 24.025 43.965 ;
		RECT	23.98 54.165 24.03 54.295 ;
		RECT	24.515 43.835 24.565 43.965 ;
		RECT	24.52 54.165 24.57 54.295 ;
		RECT	25.055 43.835 25.105 43.965 ;
		RECT	25.06 54.165 25.11 54.295 ;
		RECT	25.595 43.835 25.645 43.965 ;
		RECT	25.6 54.165 25.65 54.295 ;
		RECT	26.135 43.835 26.185 43.965 ;
		RECT	26.14 54.165 26.19 54.295 ;
		RECT	26.675 43.835 26.725 43.965 ;
		RECT	26.68 54.165 26.73 54.295 ;
		RECT	27.215 43.835 27.265 43.965 ;
		RECT	27.22 54.165 27.27 54.295 ;
		RECT	27.755 43.835 27.805 43.965 ;
		RECT	27.76 54.165 27.81 54.295 ;
		RECT	28.295 43.835 28.345 43.965 ;
		RECT	28.3 54.165 28.35 54.295 ;
		RECT	28.835 43.835 28.885 43.965 ;
		RECT	28.84 54.165 28.89 54.295 ;
		RECT	29.375 43.835 29.425 43.965 ;
		RECT	29.38 54.165 29.43 54.295 ;
		RECT	29.915 43.835 29.965 43.965 ;
		RECT	29.92 54.165 29.97 54.295 ;
		RECT	30.455 43.835 30.505 43.965 ;
		RECT	30.46 54.165 30.51 54.295 ;
		RECT	30.995 43.835 31.045 43.965 ;
		RECT	31 54.165 31.05 54.295 ;
		RECT	31.535 43.835 31.585 43.965 ;
		RECT	31.54 54.165 31.59 54.295 ;
		RECT	32.075 43.835 32.125 43.965 ;
		RECT	32.08 54.165 32.13 54.295 ;
		RECT	32.615 43.835 32.665 43.965 ;
		RECT	32.62 54.165 32.67 54.295 ;
		RECT	33.155 43.835 33.205 43.965 ;
		RECT	33.16 54.165 33.21 54.295 ;
		RECT	33.695 43.835 33.745 43.965 ;
		RECT	33.7 54.165 33.75 54.295 ;
		RECT	34.235 43.835 34.285 43.965 ;
		RECT	34.24 54.165 34.29 54.295 ;
		RECT	34.775 43.835 34.825 43.965 ;
		RECT	34.78 54.165 34.83 54.295 ;
		RECT	35.315 43.835 35.365 43.965 ;
		RECT	35.32 54.165 35.37 54.295 ;
		RECT	35.855 43.835 35.905 43.965 ;
		RECT	35.86 54.165 35.91 54.295 ;
		RECT	36.395 43.835 36.445 43.965 ;
		RECT	36.4 54.165 36.45 54.295 ;
		RECT	36.935 43.835 36.985 43.965 ;
		RECT	36.94 54.165 36.99 54.295 ;
		RECT	37.475 43.835 37.525 43.965 ;
		RECT	37.48 54.165 37.53 54.295 ;
		RECT	38.015 43.835 38.065 43.965 ;
		RECT	38.02 54.165 38.07 54.295 ;
		RECT	38.555 43.835 38.605 43.965 ;
		RECT	38.56 54.165 38.61 54.295 ;
		RECT	39.095 43.835 39.145 43.965 ;
		RECT	39.1 54.165 39.15 54.295 ;
		RECT	39.635 43.835 39.685 43.965 ;
		RECT	39.64 54.165 39.69 54.295 ;
		RECT	40.175 43.835 40.225 43.965 ;
		RECT	40.18 54.165 40.23 54.295 ;
		RECT	40.715 43.835 40.765 43.965 ;
		RECT	40.72 54.165 40.77 54.295 ;
		RECT	41.255 43.835 41.305 43.965 ;
		RECT	41.26 54.165 41.31 54.295 ;
		RECT	41.795 43.835 41.845 43.965 ;
		RECT	41.8 54.165 41.85 54.295 ;
		RECT	42.335 43.835 42.385 43.965 ;
		RECT	42.34 54.165 42.39 54.295 ;
		RECT	42.875 43.835 42.925 43.965 ;
		RECT	42.88 54.165 42.93 54.295 ;
		RECT	43.415 43.835 43.465 43.965 ;
		RECT	43.42 54.165 43.47 54.295 ;
		RECT	43.955 43.835 44.005 43.965 ;
		RECT	43.96 54.165 44.01 54.295 ;
		RECT	44.495 43.835 44.545 43.965 ;
		RECT	44.5 54.165 44.55 54.295 ;
		RECT	45.035 43.835 45.085 43.965 ;
		RECT	45.04 54.165 45.09 54.295 ;
		RECT	45.575 43.835 45.625 43.965 ;
		RECT	45.58 54.165 45.63 54.295 ;
		RECT	46.115 43.835 46.165 43.965 ;
		RECT	46.12 54.165 46.17 54.295 ;
		RECT	46.655 43.835 46.705 43.965 ;
		RECT	46.66 54.165 46.71 54.295 ;
		RECT	47.195 43.835 47.245 43.965 ;
		RECT	47.2 54.165 47.25 54.295 ;
		RECT	47.735 43.835 47.785 43.965 ;
		RECT	47.74 54.165 47.79 54.295 ;
		RECT	48.275 43.835 48.325 43.965 ;
		RECT	48.28 54.165 48.33 54.295 ;
		RECT	48.815 43.835 48.865 43.965 ;
		RECT	48.82 54.165 48.87 54.295 ;
		RECT	49.355 43.835 49.405 43.965 ;
		RECT	49.36 54.165 49.41 54.295 ;
		RECT	14.965 29.54 15.015 29.59 ;
		RECT	15.335 29.565 15.385 29.695 ;
		RECT	15.875 29.565 15.925 29.695 ;
		RECT	16.415 29.565 16.465 29.695 ;
		RECT	16.955 29.565 17.005 29.695 ;
		RECT	17.495 29.565 17.545 29.695 ;
		RECT	18.035 29.565 18.085 29.695 ;
		RECT	18.575 29.565 18.625 29.695 ;
		RECT	19.115 29.565 19.165 29.695 ;
		RECT	19.655 29.565 19.705 29.695 ;
		RECT	20.195 29.565 20.245 29.695 ;
		RECT	20.735 29.565 20.785 29.695 ;
		RECT	21.275 29.565 21.325 29.695 ;
		RECT	21.815 29.565 21.865 29.695 ;
		RECT	22.355 29.565 22.405 29.695 ;
		RECT	22.895 29.565 22.945 29.695 ;
		RECT	23.435 29.565 23.485 29.695 ;
		RECT	14.965 29.67 15.015 29.72 ;
		RECT	14.565 30.34 14.615 30.39 ;
		RECT	14.965 30.545 15.015 30.675 ;
		RECT	15.335 31.04 15.385 31.17 ;
		RECT	15.875 31.04 15.925 31.17 ;
		RECT	16.415 31.04 16.465 31.17 ;
		RECT	16.955 31.04 17.005 31.17 ;
		RECT	17.495 31.04 17.545 31.17 ;
		RECT	18.035 31.04 18.085 31.17 ;
		RECT	18.575 31.04 18.625 31.17 ;
		RECT	19.115 31.04 19.165 31.17 ;
		RECT	19.655 31.04 19.705 31.17 ;
		RECT	20.195 31.04 20.245 31.17 ;
		RECT	20.735 31.04 20.785 31.17 ;
		RECT	21.275 31.04 21.325 31.17 ;
		RECT	21.815 31.04 21.865 31.17 ;
		RECT	22.355 31.04 22.405 31.17 ;
		RECT	22.895 31.04 22.945 31.17 ;
		RECT	23.435 31.04 23.485 31.17 ;
		RECT	14.565 31.32 14.615 31.37 ;
		RECT	14.99 31.515 15.04 31.645 ;
		RECT	14.865 31.79 14.915 31.92 ;
		RECT	15.335 31.79 15.385 31.92 ;
		RECT	15.875 31.79 15.925 31.92 ;
		RECT	16.415 31.79 16.465 31.92 ;
		RECT	16.955 31.79 17.005 31.92 ;
		RECT	17.495 31.79 17.545 31.92 ;
		RECT	18.035 31.79 18.085 31.92 ;
		RECT	18.575 31.79 18.625 31.92 ;
		RECT	19.115 31.79 19.165 31.92 ;
		RECT	19.655 31.79 19.705 31.92 ;
		RECT	20.195 31.79 20.245 31.92 ;
		RECT	20.735 31.79 20.785 31.92 ;
		RECT	21.275 31.79 21.325 31.92 ;
		RECT	21.815 31.79 21.865 31.92 ;
		RECT	22.355 31.79 22.405 31.92 ;
		RECT	22.895 31.79 22.945 31.92 ;
		RECT	23.435 31.79 23.485 31.92 ;
		RECT	14.565 32.985 14.615 33.17 ;
		RECT	14.565 33.99 14.615 34.12 ;
		RECT	14.745 34.485 14.795 34.615 ;
		RECT	14.99 35.47 15.04 35.6 ;
		RECT	14.745 36.455 14.795 36.585 ;
		RECT	14.565 36.92 14.615 37.1 ;
		RECT	14.99 39.38 15.04 39.56 ;
		RECT	14.565 40.855 14.615 41.035 ;
		RECT	14.73 41.4 14.78 41.53 ;
		RECT	14.565 41.84 14.615 42.02 ;
		RECT	14.73 42.355 14.78 42.485 ;
		RECT	14.99 43.315 15.04 43.495 ;
		RECT	14.565 44.79 14.615 44.97 ;
		RECT	13.8 45.785 13.85 45.915 ;
		RECT	14.865 46.095 14.915 46.225 ;
		RECT	15.335 46.095 15.385 46.225 ;
		RECT	15.875 46.095 15.925 46.225 ;
		RECT	16.415 46.095 16.465 46.225 ;
		RECT	16.955 46.095 17.005 46.225 ;
		RECT	17.495 46.095 17.545 46.225 ;
		RECT	18.035 46.095 18.085 46.225 ;
		RECT	18.575 46.095 18.625 46.225 ;
		RECT	19.115 46.095 19.165 46.225 ;
		RECT	19.655 46.095 19.705 46.225 ;
		RECT	20.195 46.095 20.245 46.225 ;
		RECT	20.735 46.095 20.785 46.225 ;
		RECT	21.275 46.095 21.325 46.225 ;
		RECT	21.815 46.095 21.865 46.225 ;
		RECT	22.355 46.095 22.405 46.225 ;
		RECT	22.895 46.095 22.945 46.225 ;
		RECT	23.435 46.095 23.485 46.225 ;
		RECT	15.335 46.41 15.385 46.54 ;
		RECT	15.875 46.41 15.925 46.54 ;
		RECT	16.415 46.41 16.465 46.54 ;
		RECT	16.955 46.41 17.005 46.54 ;
		RECT	17.495 46.41 17.545 46.54 ;
		RECT	18.035 46.41 18.085 46.54 ;
		RECT	18.575 46.41 18.625 46.54 ;
		RECT	19.115 46.41 19.165 46.54 ;
		RECT	19.655 46.41 19.705 46.54 ;
		RECT	20.195 46.41 20.245 46.54 ;
		RECT	20.735 46.41 20.785 46.54 ;
		RECT	21.275 46.41 21.325 46.54 ;
		RECT	21.815 46.41 21.865 46.54 ;
		RECT	22.355 46.41 22.405 46.54 ;
		RECT	22.895 46.41 22.945 46.54 ;
		RECT	23.435 46.41 23.485 46.54 ;
		RECT	14.565 47.07 14.615 47.12 ;
		RECT	14.965 47.275 15.015 47.405 ;
		RECT	14.565 47.565 14.615 47.615 ;
		RECT	15.335 48.26 15.385 48.39 ;
		RECT	15.875 48.26 15.925 48.39 ;
		RECT	16.415 48.26 16.465 48.39 ;
		RECT	16.955 48.26 17.005 48.39 ;
		RECT	17.495 48.26 17.545 48.39 ;
		RECT	18.035 48.26 18.085 48.39 ;
		RECT	18.575 48.26 18.625 48.39 ;
		RECT	19.115 48.26 19.165 48.39 ;
		RECT	19.655 48.26 19.705 48.39 ;
		RECT	20.195 48.26 20.245 48.39 ;
		RECT	20.735 48.26 20.785 48.39 ;
		RECT	21.275 48.26 21.325 48.39 ;
		RECT	21.815 48.26 21.865 48.39 ;
		RECT	22.355 48.26 22.405 48.39 ;
		RECT	22.895 48.26 22.945 48.39 ;
		RECT	23.435 48.26 23.485 48.39 ;
		RECT	14.565 48.725 14.615 48.905 ;
		RECT	14.565 49.22 14.615 49.4 ;
		RECT	15.335 49.735 15.385 49.865 ;
		RECT	15.875 49.735 15.925 49.865 ;
		RECT	16.415 49.735 16.465 49.865 ;
		RECT	16.955 49.735 17.005 49.865 ;
		RECT	17.495 49.735 17.545 49.865 ;
		RECT	18.035 49.735 18.085 49.865 ;
		RECT	18.575 49.735 18.625 49.865 ;
		RECT	19.115 49.735 19.165 49.865 ;
		RECT	19.655 49.735 19.705 49.865 ;
		RECT	20.195 49.735 20.245 49.865 ;
		RECT	20.735 49.735 20.785 49.865 ;
		RECT	21.275 49.735 21.325 49.865 ;
		RECT	21.815 49.735 21.865 49.865 ;
		RECT	22.355 49.735 22.405 49.865 ;
		RECT	22.895 49.735 22.945 49.865 ;
		RECT	23.435 49.735 23.485 49.865 ;
		RECT	14.565 50.515 14.615 50.565 ;
		RECT	14.965 50.72 15.015 50.85 ;
		RECT	14.565 51.005 14.615 51.055 ;
		RECT	15.335 51.525 15.385 51.655 ;
		RECT	15.875 51.525 15.925 51.655 ;
		RECT	16.415 51.525 16.465 51.655 ;
		RECT	16.955 51.525 17.005 51.655 ;
		RECT	17.495 51.525 17.545 51.655 ;
		RECT	18.035 51.525 18.085 51.655 ;
		RECT	18.575 51.525 18.625 51.655 ;
		RECT	19.115 51.525 19.165 51.655 ;
		RECT	19.655 51.525 19.705 51.655 ;
		RECT	20.195 51.525 20.245 51.655 ;
		RECT	20.735 51.525 20.785 51.655 ;
		RECT	21.275 51.525 21.325 51.655 ;
		RECT	21.815 51.525 21.865 51.655 ;
		RECT	22.355 51.525 22.405 51.655 ;
		RECT	22.895 51.525 22.945 51.655 ;
		RECT	23.435 51.525 23.485 51.655 ;
		RECT	14.865 51.87 14.915 52 ;
		RECT	15.335 51.87 15.385 52 ;
		RECT	15.875 51.87 15.925 52 ;
		RECT	16.415 51.87 16.465 52 ;
		RECT	16.955 51.87 17.005 52 ;
		RECT	17.495 51.87 17.545 52 ;
		RECT	18.035 51.87 18.085 52 ;
		RECT	18.575 51.87 18.625 52 ;
		RECT	19.115 51.87 19.165 52 ;
		RECT	19.655 51.87 19.705 52 ;
		RECT	20.195 51.87 20.245 52 ;
		RECT	20.735 51.87 20.785 52 ;
		RECT	21.275 51.87 21.325 52 ;
		RECT	21.815 51.87 21.865 52 ;
		RECT	22.355 51.87 22.405 52 ;
		RECT	22.895 51.87 22.945 52 ;
		RECT	23.435 51.87 23.485 52 ;
		RECT	13.8 52.21 13.85 52.34 ;
		RECT	14.565 53.18 14.615 53.31 ;
		RECT	14.735 53.695 14.785 53.825 ;
		RECT	14.99 54.63 15.04 54.81 ;
		RECT	14.735 55.64 14.785 55.77 ;
		RECT	14.565 56.11 14.615 56.29 ;
		RECT	14.735 56.625 14.785 56.755 ;
		RECT	14.565 57.09 14.615 57.27 ;
		RECT	14.99 58.57 15.04 58.75 ;
		RECT	14.565 61.03 14.615 61.21 ;
		RECT	14.74 61.545 14.79 61.675 ;
		RECT	14.74 62.32 14.79 62.37 ;
		RECT	14.99 62.505 15.04 62.685 ;
		RECT	14.745 63.515 14.795 63.645 ;
		RECT	14.565 64.005 14.615 64.135 ;
		RECT	14.565 64.93 14.615 65.11 ;
		RECT	14.865 66.21 14.915 66.34 ;
		RECT	15.335 66.21 15.385 66.34 ;
		RECT	15.875 66.21 15.925 66.34 ;
		RECT	16.415 66.21 16.465 66.34 ;
		RECT	16.955 66.21 17.005 66.34 ;
		RECT	17.495 66.21 17.545 66.34 ;
		RECT	18.035 66.21 18.085 66.34 ;
		RECT	18.575 66.21 18.625 66.34 ;
		RECT	19.115 66.21 19.165 66.34 ;
		RECT	19.655 66.21 19.705 66.34 ;
		RECT	20.195 66.21 20.245 66.34 ;
		RECT	20.735 66.21 20.785 66.34 ;
		RECT	21.275 66.21 21.325 66.34 ;
		RECT	21.815 66.21 21.865 66.34 ;
		RECT	22.355 66.21 22.405 66.34 ;
		RECT	22.895 66.21 22.945 66.34 ;
		RECT	23.435 66.21 23.485 66.34 ;
		RECT	14.99 66.48 15.04 66.61 ;
		RECT	14.565 66.755 14.615 66.805 ;
		RECT	15.335 66.955 15.385 67.085 ;
		RECT	15.875 66.955 15.925 67.085 ;
		RECT	16.415 66.955 16.465 67.085 ;
		RECT	16.955 66.955 17.005 67.085 ;
		RECT	17.495 66.955 17.545 67.085 ;
		RECT	18.035 66.955 18.085 67.085 ;
		RECT	18.575 66.955 18.625 67.085 ;
		RECT	19.115 66.955 19.165 67.085 ;
		RECT	19.655 66.955 19.705 67.085 ;
		RECT	20.195 66.955 20.245 67.085 ;
		RECT	20.735 66.955 20.785 67.085 ;
		RECT	21.275 66.955 21.325 67.085 ;
		RECT	21.815 66.955 21.865 67.085 ;
		RECT	22.355 66.955 22.405 67.085 ;
		RECT	22.895 66.955 22.945 67.085 ;
		RECT	23.435 66.955 23.485 67.085 ;
		RECT	14.965 67.45 15.015 67.58 ;
		RECT	14.565 67.735 14.615 67.785 ;
		RECT	14.965 68.435 15.015 68.565 ;
		RECT	15.335 68.435 15.385 68.565 ;
		RECT	15.875 68.435 15.925 68.565 ;
		RECT	16.415 68.435 16.465 68.565 ;
		RECT	16.955 68.435 17.005 68.565 ;
		RECT	17.495 68.435 17.545 68.565 ;
		RECT	18.035 68.435 18.085 68.565 ;
		RECT	18.575 68.435 18.625 68.565 ;
		RECT	19.115 68.435 19.165 68.565 ;
		RECT	19.655 68.435 19.705 68.565 ;
		RECT	20.195 68.435 20.245 68.565 ;
		RECT	20.735 68.435 20.785 68.565 ;
		RECT	21.275 68.435 21.325 68.565 ;
		RECT	21.815 68.435 21.865 68.565 ;
		RECT	22.355 68.435 22.405 68.565 ;
		RECT	22.895 68.435 22.945 68.565 ;
		RECT	23.435 68.435 23.485 68.565 ;
		RECT	23.975 29.565 24.025 29.695 ;
		RECT	23.975 31.04 24.025 31.17 ;
		RECT	23.975 31.79 24.025 31.92 ;
		RECT	23.975 33.785 24.025 33.835 ;
		RECT	23.975 34.985 24.025 35.115 ;
		RECT	23.975 35.96 24.025 36.09 ;
		RECT	23.975 37.435 24.025 37.565 ;
		RECT	23.975 38.42 24.025 38.55 ;
		RECT	23.975 39.9 24.025 40.03 ;
		RECT	23.975 40.39 24.025 40.52 ;
		RECT	23.975 42.85 24.025 42.98 ;
		RECT	23.975 44.31 24.025 44.44 ;
		RECT	23.975 46.095 24.025 46.225 ;
		RECT	23.975 46.41 24.025 46.54 ;
		RECT	23.975 48.26 24.025 48.39 ;
		RECT	23.975 49.735 24.025 49.865 ;
		RECT	23.975 51.525 24.025 51.655 ;
		RECT	23.975 51.87 24.025 52 ;
		RECT	23.98 53.675 24.03 53.805 ;
		RECT	23.98 55.15 24.03 55.28 ;
		RECT	23.98 58.1 24.03 58.23 ;
		RECT	23.98 59.575 24.03 59.705 ;
		RECT	23.98 60.56 24.03 60.69 ;
		RECT	23.98 62.035 24.03 62.165 ;
		RECT	23.975 62.32 24.025 62.37 ;
		RECT	23.98 63.02 24.03 63.15 ;
		RECT	23.975 66.21 24.025 66.34 ;
		RECT	23.975 66.955 24.025 67.085 ;
		RECT	23.975 68.435 24.025 68.565 ;
		RECT	24.515 29.565 24.565 29.695 ;
		RECT	24.515 31.04 24.565 31.17 ;
		RECT	24.515 31.79 24.565 31.92 ;
		RECT	24.515 33.785 24.565 33.835 ;
		RECT	24.515 34.985 24.565 35.115 ;
		RECT	24.515 35.96 24.565 36.09 ;
		RECT	24.515 37.435 24.565 37.565 ;
		RECT	24.515 38.42 24.565 38.55 ;
		RECT	24.515 39.9 24.565 40.03 ;
		RECT	24.515 40.39 24.565 40.52 ;
		RECT	24.515 42.85 24.565 42.98 ;
		RECT	24.515 44.31 24.565 44.44 ;
		RECT	24.515 46.095 24.565 46.225 ;
		RECT	24.515 46.41 24.565 46.54 ;
		RECT	24.515 48.26 24.565 48.39 ;
		RECT	24.515 49.735 24.565 49.865 ;
		RECT	24.515 51.525 24.565 51.655 ;
		RECT	24.515 51.87 24.565 52 ;
		RECT	24.52 53.675 24.57 53.805 ;
		RECT	24.52 55.15 24.57 55.28 ;
		RECT	24.52 58.1 24.57 58.23 ;
		RECT	24.52 59.575 24.57 59.705 ;
		RECT	24.52 60.56 24.57 60.69 ;
		RECT	24.52 62.035 24.57 62.165 ;
		RECT	24.515 62.32 24.565 62.37 ;
		RECT	24.52 63.02 24.57 63.15 ;
		RECT	24.515 66.21 24.565 66.34 ;
		RECT	24.515 66.955 24.565 67.085 ;
		RECT	24.515 68.435 24.565 68.565 ;
		RECT	25.055 29.565 25.105 29.695 ;
		RECT	25.055 31.04 25.105 31.17 ;
		RECT	25.055 31.79 25.105 31.92 ;
		RECT	25.055 33.785 25.105 33.835 ;
		RECT	25.055 34.985 25.105 35.115 ;
		RECT	25.055 35.96 25.105 36.09 ;
		RECT	25.055 37.435 25.105 37.565 ;
		RECT	25.055 38.42 25.105 38.55 ;
		RECT	25.055 39.9 25.105 40.03 ;
		RECT	25.055 40.39 25.105 40.52 ;
		RECT	25.055 42.85 25.105 42.98 ;
		RECT	25.055 44.31 25.105 44.44 ;
		RECT	25.055 46.095 25.105 46.225 ;
		RECT	25.055 46.41 25.105 46.54 ;
		RECT	25.055 48.26 25.105 48.39 ;
		RECT	25.055 49.735 25.105 49.865 ;
		RECT	25.055 51.525 25.105 51.655 ;
		RECT	25.055 51.87 25.105 52 ;
		RECT	25.06 53.675 25.11 53.805 ;
		RECT	25.06 55.15 25.11 55.28 ;
		RECT	25.06 58.1 25.11 58.23 ;
		RECT	25.06 59.575 25.11 59.705 ;
		RECT	25.06 60.56 25.11 60.69 ;
		RECT	25.06 62.035 25.11 62.165 ;
		RECT	25.055 62.32 25.105 62.37 ;
		RECT	25.06 63.02 25.11 63.15 ;
		RECT	25.055 66.21 25.105 66.34 ;
		RECT	25.055 66.955 25.105 67.085 ;
		RECT	25.055 68.435 25.105 68.565 ;
		RECT	25.595 29.565 25.645 29.695 ;
		RECT	25.595 31.04 25.645 31.17 ;
		RECT	25.595 31.79 25.645 31.92 ;
		RECT	25.595 33.785 25.645 33.835 ;
		RECT	25.595 34.985 25.645 35.115 ;
		RECT	25.595 35.96 25.645 36.09 ;
		RECT	25.595 37.435 25.645 37.565 ;
		RECT	25.595 38.42 25.645 38.55 ;
		RECT	25.595 39.9 25.645 40.03 ;
		RECT	25.595 40.39 25.645 40.52 ;
		RECT	25.595 42.85 25.645 42.98 ;
		RECT	25.595 44.31 25.645 44.44 ;
		RECT	25.595 46.095 25.645 46.225 ;
		RECT	25.595 46.41 25.645 46.54 ;
		RECT	25.595 48.26 25.645 48.39 ;
		RECT	25.595 49.735 25.645 49.865 ;
		RECT	25.595 51.525 25.645 51.655 ;
		RECT	25.595 51.87 25.645 52 ;
		RECT	25.6 53.675 25.65 53.805 ;
		RECT	25.6 55.15 25.65 55.28 ;
		RECT	25.6 58.1 25.65 58.23 ;
		RECT	25.6 59.575 25.65 59.705 ;
		RECT	25.6 60.56 25.65 60.69 ;
		RECT	25.6 62.035 25.65 62.165 ;
		RECT	25.595 62.32 25.645 62.37 ;
		RECT	25.6 63.02 25.65 63.15 ;
		RECT	25.595 66.21 25.645 66.34 ;
		RECT	25.595 66.955 25.645 67.085 ;
		RECT	25.595 68.435 25.645 68.565 ;
		RECT	26.135 29.565 26.185 29.695 ;
		RECT	26.135 31.04 26.185 31.17 ;
		RECT	26.135 31.79 26.185 31.92 ;
		RECT	26.135 33.785 26.185 33.835 ;
		RECT	26.135 34.985 26.185 35.115 ;
		RECT	26.135 35.96 26.185 36.09 ;
		RECT	26.135 37.435 26.185 37.565 ;
		RECT	26.135 38.42 26.185 38.55 ;
		RECT	26.135 39.9 26.185 40.03 ;
		RECT	26.135 40.39 26.185 40.52 ;
		RECT	26.135 42.85 26.185 42.98 ;
		RECT	26.135 44.31 26.185 44.44 ;
		RECT	26.135 46.095 26.185 46.225 ;
		RECT	26.135 46.41 26.185 46.54 ;
		RECT	26.135 48.26 26.185 48.39 ;
		RECT	26.135 49.735 26.185 49.865 ;
		RECT	26.135 51.525 26.185 51.655 ;
		RECT	26.135 51.87 26.185 52 ;
		RECT	26.14 53.675 26.19 53.805 ;
		RECT	26.14 55.15 26.19 55.28 ;
		RECT	26.14 58.1 26.19 58.23 ;
		RECT	26.14 59.575 26.19 59.705 ;
		RECT	26.14 60.56 26.19 60.69 ;
		RECT	26.14 62.035 26.19 62.165 ;
		RECT	26.135 62.32 26.185 62.37 ;
		RECT	26.14 63.02 26.19 63.15 ;
		RECT	26.135 66.21 26.185 66.34 ;
		RECT	26.135 66.955 26.185 67.085 ;
		RECT	26.135 68.435 26.185 68.565 ;
		RECT	26.675 29.565 26.725 29.695 ;
		RECT	26.675 31.04 26.725 31.17 ;
		RECT	26.675 31.79 26.725 31.92 ;
		RECT	26.675 33.785 26.725 33.835 ;
		RECT	26.675 34.985 26.725 35.115 ;
		RECT	26.675 35.96 26.725 36.09 ;
		RECT	26.675 37.435 26.725 37.565 ;
		RECT	26.675 38.42 26.725 38.55 ;
		RECT	26.675 39.9 26.725 40.03 ;
		RECT	26.675 40.39 26.725 40.52 ;
		RECT	26.675 42.85 26.725 42.98 ;
		RECT	26.675 44.31 26.725 44.44 ;
		RECT	26.675 46.095 26.725 46.225 ;
		RECT	26.675 46.41 26.725 46.54 ;
		RECT	26.675 48.26 26.725 48.39 ;
		RECT	26.675 49.735 26.725 49.865 ;
		RECT	26.675 51.525 26.725 51.655 ;
		RECT	26.675 51.87 26.725 52 ;
		RECT	26.68 53.675 26.73 53.805 ;
		RECT	26.68 55.15 26.73 55.28 ;
		RECT	26.68 58.1 26.73 58.23 ;
		RECT	26.68 59.575 26.73 59.705 ;
		RECT	26.68 60.56 26.73 60.69 ;
		RECT	26.68 62.035 26.73 62.165 ;
		RECT	26.675 62.32 26.725 62.37 ;
		RECT	26.68 63.02 26.73 63.15 ;
		RECT	26.675 66.21 26.725 66.34 ;
		RECT	26.675 66.955 26.725 67.085 ;
		RECT	26.675 68.435 26.725 68.565 ;
		RECT	27.215 29.565 27.265 29.695 ;
		RECT	27.215 31.04 27.265 31.17 ;
		RECT	27.215 31.79 27.265 31.92 ;
		RECT	27.215 33.785 27.265 33.835 ;
		RECT	27.215 34.985 27.265 35.115 ;
		RECT	27.215 35.96 27.265 36.09 ;
		RECT	27.215 37.435 27.265 37.565 ;
		RECT	27.215 38.42 27.265 38.55 ;
		RECT	27.215 39.9 27.265 40.03 ;
		RECT	27.215 40.39 27.265 40.52 ;
		RECT	27.215 42.85 27.265 42.98 ;
		RECT	27.215 44.31 27.265 44.44 ;
		RECT	27.215 46.095 27.265 46.225 ;
		RECT	27.215 46.41 27.265 46.54 ;
		RECT	27.215 48.26 27.265 48.39 ;
		RECT	27.215 49.735 27.265 49.865 ;
		RECT	27.215 51.525 27.265 51.655 ;
		RECT	27.215 51.87 27.265 52 ;
		RECT	27.22 53.675 27.27 53.805 ;
		RECT	27.22 55.15 27.27 55.28 ;
		RECT	27.22 58.1 27.27 58.23 ;
		RECT	27.22 59.575 27.27 59.705 ;
		RECT	27.22 60.56 27.27 60.69 ;
		RECT	27.22 62.035 27.27 62.165 ;
		RECT	27.215 62.32 27.265 62.37 ;
		RECT	27.22 63.02 27.27 63.15 ;
		RECT	27.215 66.21 27.265 66.34 ;
		RECT	27.215 66.955 27.265 67.085 ;
		RECT	27.215 68.435 27.265 68.565 ;
		RECT	27.755 29.565 27.805 29.695 ;
		RECT	27.755 31.04 27.805 31.17 ;
		RECT	27.755 31.79 27.805 31.92 ;
		RECT	27.755 33.785 27.805 33.835 ;
		RECT	27.755 34.985 27.805 35.115 ;
		RECT	27.755 35.96 27.805 36.09 ;
		RECT	27.755 37.435 27.805 37.565 ;
		RECT	27.755 38.42 27.805 38.55 ;
		RECT	27.755 39.9 27.805 40.03 ;
		RECT	27.755 40.39 27.805 40.52 ;
		RECT	27.755 42.85 27.805 42.98 ;
		RECT	27.755 44.31 27.805 44.44 ;
		RECT	27.755 46.095 27.805 46.225 ;
		RECT	27.755 46.41 27.805 46.54 ;
		RECT	27.755 48.26 27.805 48.39 ;
		RECT	27.755 49.735 27.805 49.865 ;
		RECT	27.755 51.525 27.805 51.655 ;
		RECT	27.755 51.87 27.805 52 ;
		RECT	27.76 53.675 27.81 53.805 ;
		RECT	27.76 55.15 27.81 55.28 ;
		RECT	27.76 58.1 27.81 58.23 ;
		RECT	27.76 59.575 27.81 59.705 ;
		RECT	27.76 60.56 27.81 60.69 ;
		RECT	27.76 62.035 27.81 62.165 ;
		RECT	27.755 62.32 27.805 62.37 ;
		RECT	27.76 63.02 27.81 63.15 ;
		RECT	27.755 66.21 27.805 66.34 ;
		RECT	27.755 66.955 27.805 67.085 ;
		RECT	27.755 68.435 27.805 68.565 ;
		RECT	28.295 29.565 28.345 29.695 ;
		RECT	28.295 31.04 28.345 31.17 ;
		RECT	28.295 31.79 28.345 31.92 ;
		RECT	28.295 33.785 28.345 33.835 ;
		RECT	28.295 34.985 28.345 35.115 ;
		RECT	28.295 35.96 28.345 36.09 ;
		RECT	28.295 37.435 28.345 37.565 ;
		RECT	28.295 38.42 28.345 38.55 ;
		RECT	28.295 39.9 28.345 40.03 ;
		RECT	28.295 40.39 28.345 40.52 ;
		RECT	28.295 42.85 28.345 42.98 ;
		RECT	28.295 44.31 28.345 44.44 ;
		RECT	28.295 46.095 28.345 46.225 ;
		RECT	28.295 46.41 28.345 46.54 ;
		RECT	28.295 48.26 28.345 48.39 ;
		RECT	28.295 49.735 28.345 49.865 ;
		RECT	28.295 51.525 28.345 51.655 ;
		RECT	28.295 51.87 28.345 52 ;
		RECT	28.3 53.675 28.35 53.805 ;
		RECT	28.3 55.15 28.35 55.28 ;
		RECT	28.3 58.1 28.35 58.23 ;
		RECT	28.3 59.575 28.35 59.705 ;
		RECT	28.3 60.56 28.35 60.69 ;
		RECT	28.3 62.035 28.35 62.165 ;
		RECT	28.295 62.32 28.345 62.37 ;
		RECT	28.3 63.02 28.35 63.15 ;
		RECT	28.295 66.21 28.345 66.34 ;
		RECT	28.295 66.955 28.345 67.085 ;
		RECT	28.295 68.435 28.345 68.565 ;
		RECT	28.835 29.565 28.885 29.695 ;
		RECT	28.835 31.04 28.885 31.17 ;
		RECT	28.835 31.79 28.885 31.92 ;
		RECT	28.835 33.785 28.885 33.835 ;
		RECT	28.835 34.985 28.885 35.115 ;
		RECT	28.835 35.96 28.885 36.09 ;
		RECT	28.835 37.435 28.885 37.565 ;
		RECT	28.835 38.42 28.885 38.55 ;
		RECT	28.835 39.9 28.885 40.03 ;
		RECT	28.835 40.39 28.885 40.52 ;
		RECT	28.835 42.85 28.885 42.98 ;
		RECT	28.835 44.31 28.885 44.44 ;
		RECT	28.835 46.095 28.885 46.225 ;
		RECT	28.835 46.41 28.885 46.54 ;
		RECT	28.835 48.26 28.885 48.39 ;
		RECT	28.835 49.735 28.885 49.865 ;
		RECT	28.835 51.525 28.885 51.655 ;
		RECT	28.835 51.87 28.885 52 ;
		RECT	28.84 53.675 28.89 53.805 ;
		RECT	28.84 55.15 28.89 55.28 ;
		RECT	28.84 58.1 28.89 58.23 ;
		RECT	28.84 59.575 28.89 59.705 ;
		RECT	28.84 60.56 28.89 60.69 ;
		RECT	28.84 62.035 28.89 62.165 ;
		RECT	28.835 62.32 28.885 62.37 ;
		RECT	28.84 63.02 28.89 63.15 ;
		RECT	28.835 66.21 28.885 66.34 ;
		RECT	28.835 66.955 28.885 67.085 ;
		RECT	28.835 68.435 28.885 68.565 ;
		RECT	29.375 29.565 29.425 29.695 ;
		RECT	29.375 31.04 29.425 31.17 ;
		RECT	29.375 31.79 29.425 31.92 ;
		RECT	29.375 33.785 29.425 33.835 ;
		RECT	29.375 34.985 29.425 35.115 ;
		RECT	29.375 35.96 29.425 36.09 ;
		RECT	29.375 37.435 29.425 37.565 ;
		RECT	29.375 38.42 29.425 38.55 ;
		RECT	29.375 39.9 29.425 40.03 ;
		RECT	29.375 40.39 29.425 40.52 ;
		RECT	29.375 42.85 29.425 42.98 ;
		RECT	29.375 44.31 29.425 44.44 ;
		RECT	29.375 46.095 29.425 46.225 ;
		RECT	29.375 46.41 29.425 46.54 ;
		RECT	29.375 48.26 29.425 48.39 ;
		RECT	29.375 49.735 29.425 49.865 ;
		RECT	29.375 51.525 29.425 51.655 ;
		RECT	29.375 51.87 29.425 52 ;
		RECT	29.38 53.675 29.43 53.805 ;
		RECT	29.38 55.15 29.43 55.28 ;
		RECT	29.38 58.1 29.43 58.23 ;
		RECT	29.38 59.575 29.43 59.705 ;
		RECT	29.38 60.56 29.43 60.69 ;
		RECT	29.38 62.035 29.43 62.165 ;
		RECT	29.375 62.32 29.425 62.37 ;
		RECT	29.38 63.02 29.43 63.15 ;
		RECT	29.375 66.21 29.425 66.34 ;
		RECT	29.375 66.955 29.425 67.085 ;
		RECT	29.375 68.435 29.425 68.565 ;
		RECT	29.915 29.565 29.965 29.695 ;
		RECT	29.915 31.04 29.965 31.17 ;
		RECT	29.915 31.79 29.965 31.92 ;
		RECT	29.915 33.785 29.965 33.835 ;
		RECT	29.915 34.985 29.965 35.115 ;
		RECT	29.915 35.96 29.965 36.09 ;
		RECT	29.915 37.435 29.965 37.565 ;
		RECT	29.915 38.42 29.965 38.55 ;
		RECT	29.915 39.9 29.965 40.03 ;
		RECT	29.915 40.39 29.965 40.52 ;
		RECT	29.915 42.85 29.965 42.98 ;
		RECT	29.915 44.31 29.965 44.44 ;
		RECT	29.915 46.095 29.965 46.225 ;
		RECT	29.915 46.41 29.965 46.54 ;
		RECT	29.915 48.26 29.965 48.39 ;
		RECT	29.915 49.735 29.965 49.865 ;
		RECT	29.915 51.525 29.965 51.655 ;
		RECT	29.915 51.87 29.965 52 ;
		RECT	29.92 53.675 29.97 53.805 ;
		RECT	29.92 55.15 29.97 55.28 ;
		RECT	29.92 58.1 29.97 58.23 ;
		RECT	29.92 59.575 29.97 59.705 ;
		RECT	29.92 60.56 29.97 60.69 ;
		RECT	29.92 62.035 29.97 62.165 ;
		RECT	29.915 62.32 29.965 62.37 ;
		RECT	29.92 63.02 29.97 63.15 ;
		RECT	29.915 66.21 29.965 66.34 ;
		RECT	29.915 66.955 29.965 67.085 ;
		RECT	29.915 68.435 29.965 68.565 ;
		RECT	30.455 29.565 30.505 29.695 ;
		RECT	30.455 31.04 30.505 31.17 ;
		RECT	30.455 31.79 30.505 31.92 ;
		RECT	30.455 33.785 30.505 33.835 ;
		RECT	30.455 34.985 30.505 35.115 ;
		RECT	30.455 35.96 30.505 36.09 ;
		RECT	30.455 37.435 30.505 37.565 ;
		RECT	30.455 38.42 30.505 38.55 ;
		RECT	30.455 39.9 30.505 40.03 ;
		RECT	30.455 40.39 30.505 40.52 ;
		RECT	30.455 42.85 30.505 42.98 ;
		RECT	30.455 44.31 30.505 44.44 ;
		RECT	30.455 46.095 30.505 46.225 ;
		RECT	30.455 46.41 30.505 46.54 ;
		RECT	30.455 48.26 30.505 48.39 ;
		RECT	30.455 49.735 30.505 49.865 ;
		RECT	30.455 51.525 30.505 51.655 ;
		RECT	30.455 51.87 30.505 52 ;
		RECT	30.46 53.675 30.51 53.805 ;
		RECT	30.46 55.15 30.51 55.28 ;
		RECT	30.46 58.1 30.51 58.23 ;
		RECT	30.46 59.575 30.51 59.705 ;
		RECT	30.46 60.56 30.51 60.69 ;
		RECT	30.46 62.035 30.51 62.165 ;
		RECT	30.455 62.32 30.505 62.37 ;
		RECT	30.46 63.02 30.51 63.15 ;
		RECT	30.455 66.21 30.505 66.34 ;
		RECT	30.455 66.955 30.505 67.085 ;
		RECT	30.455 68.435 30.505 68.565 ;
		RECT	30.995 29.565 31.045 29.695 ;
		RECT	30.995 31.04 31.045 31.17 ;
		RECT	30.995 31.79 31.045 31.92 ;
		RECT	30.995 33.785 31.045 33.835 ;
		RECT	30.995 34.985 31.045 35.115 ;
		RECT	30.995 35.96 31.045 36.09 ;
		RECT	30.995 37.435 31.045 37.565 ;
		RECT	30.995 38.42 31.045 38.55 ;
		RECT	30.995 39.9 31.045 40.03 ;
		RECT	30.995 40.39 31.045 40.52 ;
		RECT	30.995 42.85 31.045 42.98 ;
		RECT	30.995 44.31 31.045 44.44 ;
		RECT	30.995 46.095 31.045 46.225 ;
		RECT	30.995 46.41 31.045 46.54 ;
		RECT	30.995 48.26 31.045 48.39 ;
		RECT	30.995 49.735 31.045 49.865 ;
		RECT	30.995 51.525 31.045 51.655 ;
		RECT	30.995 51.87 31.045 52 ;
		RECT	31 53.675 31.05 53.805 ;
		RECT	31 55.15 31.05 55.28 ;
		RECT	31 58.1 31.05 58.23 ;
		RECT	31 59.575 31.05 59.705 ;
		RECT	31 60.56 31.05 60.69 ;
		RECT	31 62.035 31.05 62.165 ;
		RECT	30.995 62.32 31.045 62.37 ;
		RECT	31 63.02 31.05 63.15 ;
		RECT	30.995 66.21 31.045 66.34 ;
		RECT	30.995 66.955 31.045 67.085 ;
		RECT	30.995 68.435 31.045 68.565 ;
		RECT	31.535 29.565 31.585 29.695 ;
		RECT	31.535 31.04 31.585 31.17 ;
		RECT	31.535 31.79 31.585 31.92 ;
		RECT	31.535 33.785 31.585 33.835 ;
		RECT	31.535 34.985 31.585 35.115 ;
		RECT	31.535 35.96 31.585 36.09 ;
		RECT	31.535 37.435 31.585 37.565 ;
		RECT	31.535 38.42 31.585 38.55 ;
		RECT	31.535 39.9 31.585 40.03 ;
		RECT	31.535 40.39 31.585 40.52 ;
		RECT	31.535 42.85 31.585 42.98 ;
		RECT	31.535 44.31 31.585 44.44 ;
		RECT	31.535 46.095 31.585 46.225 ;
		RECT	31.535 46.41 31.585 46.54 ;
		RECT	31.535 48.26 31.585 48.39 ;
		RECT	31.535 49.735 31.585 49.865 ;
		RECT	31.535 51.525 31.585 51.655 ;
		RECT	31.535 51.87 31.585 52 ;
		RECT	31.54 53.675 31.59 53.805 ;
		RECT	31.54 55.15 31.59 55.28 ;
		RECT	31.54 58.1 31.59 58.23 ;
		RECT	31.54 59.575 31.59 59.705 ;
		RECT	31.54 60.56 31.59 60.69 ;
		RECT	31.54 62.035 31.59 62.165 ;
		RECT	31.535 62.32 31.585 62.37 ;
		RECT	31.54 63.02 31.59 63.15 ;
		RECT	31.535 66.21 31.585 66.34 ;
		RECT	31.535 66.955 31.585 67.085 ;
		RECT	31.535 68.435 31.585 68.565 ;
		RECT	32.075 29.565 32.125 29.695 ;
		RECT	32.075 31.04 32.125 31.17 ;
		RECT	32.075 31.79 32.125 31.92 ;
		RECT	32.075 33.785 32.125 33.835 ;
		RECT	32.075 34.985 32.125 35.115 ;
		RECT	32.075 35.96 32.125 36.09 ;
		RECT	32.075 37.435 32.125 37.565 ;
		RECT	32.075 38.42 32.125 38.55 ;
		RECT	32.075 39.9 32.125 40.03 ;
		RECT	32.075 40.39 32.125 40.52 ;
		RECT	32.075 42.85 32.125 42.98 ;
		RECT	32.075 44.31 32.125 44.44 ;
		RECT	32.075 46.095 32.125 46.225 ;
		RECT	32.075 46.41 32.125 46.54 ;
		RECT	32.075 48.26 32.125 48.39 ;
		RECT	32.075 49.735 32.125 49.865 ;
		RECT	32.075 51.525 32.125 51.655 ;
		RECT	32.075 51.87 32.125 52 ;
		RECT	32.08 53.675 32.13 53.805 ;
		RECT	32.08 55.15 32.13 55.28 ;
		RECT	32.08 58.1 32.13 58.23 ;
		RECT	32.08 59.575 32.13 59.705 ;
		RECT	32.08 60.56 32.13 60.69 ;
		RECT	32.08 62.035 32.13 62.165 ;
		RECT	32.075 62.32 32.125 62.37 ;
		RECT	32.08 63.02 32.13 63.15 ;
		RECT	32.075 66.21 32.125 66.34 ;
		RECT	32.075 66.955 32.125 67.085 ;
		RECT	32.075 68.435 32.125 68.565 ;
		RECT	32.615 29.565 32.665 29.695 ;
		RECT	32.615 31.04 32.665 31.17 ;
		RECT	32.615 31.79 32.665 31.92 ;
		RECT	32.615 33.785 32.665 33.835 ;
		RECT	32.615 34.985 32.665 35.115 ;
		RECT	32.615 35.96 32.665 36.09 ;
		RECT	32.615 37.435 32.665 37.565 ;
		RECT	32.615 38.42 32.665 38.55 ;
		RECT	32.615 39.9 32.665 40.03 ;
		RECT	32.615 40.39 32.665 40.52 ;
		RECT	32.615 42.85 32.665 42.98 ;
		RECT	32.615 44.31 32.665 44.44 ;
		RECT	32.615 46.095 32.665 46.225 ;
		RECT	32.615 46.41 32.665 46.54 ;
		RECT	32.615 48.26 32.665 48.39 ;
		RECT	32.615 49.735 32.665 49.865 ;
		RECT	32.615 51.525 32.665 51.655 ;
		RECT	32.615 51.87 32.665 52 ;
		RECT	32.62 53.675 32.67 53.805 ;
		RECT	32.62 55.15 32.67 55.28 ;
		RECT	32.62 58.1 32.67 58.23 ;
		RECT	32.62 59.575 32.67 59.705 ;
		RECT	32.62 60.56 32.67 60.69 ;
		RECT	32.62 62.035 32.67 62.165 ;
		RECT	32.615 62.32 32.665 62.37 ;
		RECT	32.62 63.02 32.67 63.15 ;
		RECT	32.615 66.21 32.665 66.34 ;
		RECT	32.615 66.955 32.665 67.085 ;
		RECT	32.615 68.435 32.665 68.565 ;
		RECT	33.155 29.565 33.205 29.695 ;
		RECT	33.155 31.04 33.205 31.17 ;
		RECT	33.155 31.79 33.205 31.92 ;
		RECT	33.155 33.785 33.205 33.835 ;
		RECT	33.155 34.985 33.205 35.115 ;
		RECT	33.155 35.96 33.205 36.09 ;
		RECT	33.155 37.435 33.205 37.565 ;
		RECT	33.155 38.42 33.205 38.55 ;
		RECT	33.155 39.9 33.205 40.03 ;
		RECT	33.155 40.39 33.205 40.52 ;
		RECT	33.155 42.85 33.205 42.98 ;
		RECT	33.155 44.31 33.205 44.44 ;
		RECT	33.155 46.095 33.205 46.225 ;
		RECT	33.155 46.41 33.205 46.54 ;
		RECT	33.155 48.26 33.205 48.39 ;
		RECT	33.155 49.735 33.205 49.865 ;
		RECT	33.155 51.525 33.205 51.655 ;
		RECT	33.155 51.87 33.205 52 ;
		RECT	33.16 53.675 33.21 53.805 ;
		RECT	33.16 55.15 33.21 55.28 ;
		RECT	33.16 58.1 33.21 58.23 ;
		RECT	33.16 59.575 33.21 59.705 ;
		RECT	33.16 60.56 33.21 60.69 ;
		RECT	33.16 62.035 33.21 62.165 ;
		RECT	33.155 62.32 33.205 62.37 ;
		RECT	33.16 63.02 33.21 63.15 ;
		RECT	33.155 66.21 33.205 66.34 ;
		RECT	33.155 66.955 33.205 67.085 ;
		RECT	33.155 68.435 33.205 68.565 ;
		RECT	33.695 29.565 33.745 29.695 ;
		RECT	33.695 31.04 33.745 31.17 ;
		RECT	33.695 31.79 33.745 31.92 ;
		RECT	33.695 33.785 33.745 33.835 ;
		RECT	33.695 34.985 33.745 35.115 ;
		RECT	33.695 35.96 33.745 36.09 ;
		RECT	33.695 37.435 33.745 37.565 ;
		RECT	33.695 38.42 33.745 38.55 ;
		RECT	33.695 39.9 33.745 40.03 ;
		RECT	33.695 40.39 33.745 40.52 ;
		RECT	33.695 42.85 33.745 42.98 ;
		RECT	33.695 44.31 33.745 44.44 ;
		RECT	33.695 46.095 33.745 46.225 ;
		RECT	33.695 46.41 33.745 46.54 ;
		RECT	33.695 48.26 33.745 48.39 ;
		RECT	33.695 49.735 33.745 49.865 ;
		RECT	33.695 51.525 33.745 51.655 ;
		RECT	33.695 51.87 33.745 52 ;
		RECT	33.7 53.675 33.75 53.805 ;
		RECT	33.7 55.15 33.75 55.28 ;
		RECT	33.7 58.1 33.75 58.23 ;
		RECT	33.7 59.575 33.75 59.705 ;
		RECT	33.7 60.56 33.75 60.69 ;
		RECT	33.7 62.035 33.75 62.165 ;
		RECT	33.695 62.32 33.745 62.37 ;
		RECT	33.7 63.02 33.75 63.15 ;
		RECT	33.695 66.21 33.745 66.34 ;
		RECT	33.695 66.955 33.745 67.085 ;
		RECT	33.695 68.435 33.745 68.565 ;
		RECT	34.235 29.565 34.285 29.695 ;
		RECT	34.235 31.04 34.285 31.17 ;
		RECT	34.235 31.79 34.285 31.92 ;
		RECT	34.235 33.785 34.285 33.835 ;
		RECT	34.235 34.985 34.285 35.115 ;
		RECT	34.235 35.96 34.285 36.09 ;
		RECT	34.235 37.435 34.285 37.565 ;
		RECT	34.235 38.42 34.285 38.55 ;
		RECT	34.235 39.9 34.285 40.03 ;
		RECT	34.235 40.39 34.285 40.52 ;
		RECT	34.235 42.85 34.285 42.98 ;
		RECT	34.235 44.31 34.285 44.44 ;
		RECT	34.235 46.095 34.285 46.225 ;
		RECT	34.235 46.41 34.285 46.54 ;
		RECT	34.235 48.26 34.285 48.39 ;
		RECT	34.235 49.735 34.285 49.865 ;
		RECT	34.235 51.525 34.285 51.655 ;
		RECT	34.235 51.87 34.285 52 ;
		RECT	34.24 53.675 34.29 53.805 ;
		RECT	34.24 55.15 34.29 55.28 ;
		RECT	34.24 58.1 34.29 58.23 ;
		RECT	34.24 59.575 34.29 59.705 ;
		RECT	34.24 60.56 34.29 60.69 ;
		RECT	34.24 62.035 34.29 62.165 ;
		RECT	34.235 62.32 34.285 62.37 ;
		RECT	34.24 63.02 34.29 63.15 ;
		RECT	34.235 66.21 34.285 66.34 ;
		RECT	34.235 66.955 34.285 67.085 ;
		RECT	34.235 68.435 34.285 68.565 ;
		RECT	34.775 29.565 34.825 29.695 ;
		RECT	34.775 31.04 34.825 31.17 ;
		RECT	34.775 31.79 34.825 31.92 ;
		RECT	34.775 33.785 34.825 33.835 ;
		RECT	34.775 34.985 34.825 35.115 ;
		RECT	34.775 35.96 34.825 36.09 ;
		RECT	34.775 37.435 34.825 37.565 ;
		RECT	34.775 38.42 34.825 38.55 ;
		RECT	34.775 39.9 34.825 40.03 ;
		RECT	34.775 40.39 34.825 40.52 ;
		RECT	34.775 42.85 34.825 42.98 ;
		RECT	34.775 44.31 34.825 44.44 ;
		RECT	34.775 46.095 34.825 46.225 ;
		RECT	34.775 46.41 34.825 46.54 ;
		RECT	34.775 48.26 34.825 48.39 ;
		RECT	34.775 49.735 34.825 49.865 ;
		RECT	34.775 51.525 34.825 51.655 ;
		RECT	34.775 51.87 34.825 52 ;
		RECT	34.78 53.675 34.83 53.805 ;
		RECT	34.78 55.15 34.83 55.28 ;
		RECT	34.78 58.1 34.83 58.23 ;
		RECT	34.78 59.575 34.83 59.705 ;
		RECT	34.78 60.56 34.83 60.69 ;
		RECT	34.78 62.035 34.83 62.165 ;
		RECT	34.775 62.32 34.825 62.37 ;
		RECT	34.78 63.02 34.83 63.15 ;
		RECT	34.775 66.21 34.825 66.34 ;
		RECT	34.775 66.955 34.825 67.085 ;
		RECT	34.775 68.435 34.825 68.565 ;
		RECT	35.315 29.565 35.365 29.695 ;
		RECT	35.315 31.04 35.365 31.17 ;
		RECT	35.315 31.79 35.365 31.92 ;
		RECT	35.315 33.785 35.365 33.835 ;
		RECT	35.315 34.985 35.365 35.115 ;
		RECT	35.315 35.96 35.365 36.09 ;
		RECT	35.315 37.435 35.365 37.565 ;
		RECT	35.315 38.42 35.365 38.55 ;
		RECT	35.315 39.9 35.365 40.03 ;
		RECT	35.315 40.39 35.365 40.52 ;
		RECT	35.315 42.85 35.365 42.98 ;
		RECT	35.315 44.31 35.365 44.44 ;
		RECT	35.315 46.095 35.365 46.225 ;
		RECT	35.315 46.41 35.365 46.54 ;
		RECT	35.315 48.26 35.365 48.39 ;
		RECT	35.315 49.735 35.365 49.865 ;
		RECT	35.315 51.525 35.365 51.655 ;
		RECT	35.315 51.87 35.365 52 ;
		RECT	35.32 53.675 35.37 53.805 ;
		RECT	35.32 55.15 35.37 55.28 ;
		RECT	35.32 58.1 35.37 58.23 ;
		RECT	35.32 59.575 35.37 59.705 ;
		RECT	35.32 60.56 35.37 60.69 ;
		RECT	35.32 62.035 35.37 62.165 ;
		RECT	35.315 62.32 35.365 62.37 ;
		RECT	35.32 63.02 35.37 63.15 ;
		RECT	35.315 66.21 35.365 66.34 ;
		RECT	35.315 66.955 35.365 67.085 ;
		RECT	35.315 68.435 35.365 68.565 ;
		RECT	35.855 29.565 35.905 29.695 ;
		RECT	35.855 31.04 35.905 31.17 ;
		RECT	35.855 31.79 35.905 31.92 ;
		RECT	35.855 33.785 35.905 33.835 ;
		RECT	35.855 34.985 35.905 35.115 ;
		RECT	35.855 35.96 35.905 36.09 ;
		RECT	35.855 37.435 35.905 37.565 ;
		RECT	35.855 38.42 35.905 38.55 ;
		RECT	35.855 39.9 35.905 40.03 ;
		RECT	35.855 40.39 35.905 40.52 ;
		RECT	35.855 42.85 35.905 42.98 ;
		RECT	35.855 44.31 35.905 44.44 ;
		RECT	35.855 46.095 35.905 46.225 ;
		RECT	35.855 46.41 35.905 46.54 ;
		RECT	35.855 48.26 35.905 48.39 ;
		RECT	35.855 49.735 35.905 49.865 ;
		RECT	35.855 51.525 35.905 51.655 ;
		RECT	35.855 51.87 35.905 52 ;
		RECT	35.86 53.675 35.91 53.805 ;
		RECT	35.86 55.15 35.91 55.28 ;
		RECT	35.86 58.1 35.91 58.23 ;
		RECT	35.86 59.575 35.91 59.705 ;
		RECT	35.86 60.56 35.91 60.69 ;
		RECT	35.86 62.035 35.91 62.165 ;
		RECT	35.855 62.32 35.905 62.37 ;
		RECT	35.86 63.02 35.91 63.15 ;
		RECT	35.855 66.21 35.905 66.34 ;
		RECT	35.855 66.955 35.905 67.085 ;
		RECT	35.855 68.435 35.905 68.565 ;
		RECT	36.395 29.565 36.445 29.695 ;
		RECT	36.395 31.04 36.445 31.17 ;
		RECT	36.395 31.79 36.445 31.92 ;
		RECT	36.395 33.785 36.445 33.835 ;
		RECT	36.395 34.985 36.445 35.115 ;
		RECT	36.395 35.96 36.445 36.09 ;
		RECT	36.395 37.435 36.445 37.565 ;
		RECT	36.395 38.42 36.445 38.55 ;
		RECT	36.395 39.9 36.445 40.03 ;
		RECT	36.395 40.39 36.445 40.52 ;
		RECT	36.395 42.85 36.445 42.98 ;
		RECT	36.395 44.31 36.445 44.44 ;
		RECT	36.395 46.095 36.445 46.225 ;
		RECT	36.395 46.41 36.445 46.54 ;
		RECT	36.395 48.26 36.445 48.39 ;
		RECT	36.395 49.735 36.445 49.865 ;
		RECT	36.395 51.525 36.445 51.655 ;
		RECT	36.395 51.87 36.445 52 ;
		RECT	36.4 53.675 36.45 53.805 ;
		RECT	36.4 55.15 36.45 55.28 ;
		RECT	36.4 58.1 36.45 58.23 ;
		RECT	36.4 59.575 36.45 59.705 ;
		RECT	36.4 60.56 36.45 60.69 ;
		RECT	36.4 62.035 36.45 62.165 ;
		RECT	36.395 62.32 36.445 62.37 ;
		RECT	36.4 63.02 36.45 63.15 ;
		RECT	36.395 66.21 36.445 66.34 ;
		RECT	36.395 66.955 36.445 67.085 ;
		RECT	36.395 68.435 36.445 68.565 ;
		RECT	36.935 29.565 36.985 29.695 ;
		RECT	36.935 31.04 36.985 31.17 ;
		RECT	36.935 31.79 36.985 31.92 ;
		RECT	36.935 33.785 36.985 33.835 ;
		RECT	36.935 34.985 36.985 35.115 ;
		RECT	36.935 35.96 36.985 36.09 ;
		RECT	36.935 37.435 36.985 37.565 ;
		RECT	36.935 38.42 36.985 38.55 ;
		RECT	36.935 39.9 36.985 40.03 ;
		RECT	36.935 40.39 36.985 40.52 ;
		RECT	36.935 42.85 36.985 42.98 ;
		RECT	36.935 44.31 36.985 44.44 ;
		RECT	36.935 46.095 36.985 46.225 ;
		RECT	36.935 46.41 36.985 46.54 ;
		RECT	36.935 48.26 36.985 48.39 ;
		RECT	36.935 49.735 36.985 49.865 ;
		RECT	36.935 51.525 36.985 51.655 ;
		RECT	36.935 51.87 36.985 52 ;
		RECT	36.94 53.675 36.99 53.805 ;
		RECT	36.94 55.15 36.99 55.28 ;
		RECT	36.94 58.1 36.99 58.23 ;
		RECT	36.94 59.575 36.99 59.705 ;
		RECT	36.94 60.56 36.99 60.69 ;
		RECT	36.94 62.035 36.99 62.165 ;
		RECT	36.935 62.32 36.985 62.37 ;
		RECT	36.94 63.02 36.99 63.15 ;
		RECT	36.935 66.21 36.985 66.34 ;
		RECT	36.935 66.955 36.985 67.085 ;
		RECT	36.935 68.435 36.985 68.565 ;
		RECT	37.475 29.565 37.525 29.695 ;
		RECT	37.475 31.04 37.525 31.17 ;
		RECT	37.475 31.79 37.525 31.92 ;
		RECT	37.475 33.785 37.525 33.835 ;
		RECT	37.475 34.985 37.525 35.115 ;
		RECT	37.475 35.96 37.525 36.09 ;
		RECT	37.475 37.435 37.525 37.565 ;
		RECT	37.475 38.42 37.525 38.55 ;
		RECT	37.475 39.9 37.525 40.03 ;
		RECT	37.475 40.39 37.525 40.52 ;
		RECT	37.475 42.85 37.525 42.98 ;
		RECT	37.475 44.31 37.525 44.44 ;
		RECT	37.475 46.095 37.525 46.225 ;
		RECT	37.475 46.41 37.525 46.54 ;
		RECT	37.475 48.26 37.525 48.39 ;
		RECT	37.475 49.735 37.525 49.865 ;
		RECT	37.475 51.525 37.525 51.655 ;
		RECT	37.475 51.87 37.525 52 ;
		RECT	37.48 53.675 37.53 53.805 ;
		RECT	37.48 55.15 37.53 55.28 ;
		RECT	37.48 58.1 37.53 58.23 ;
		RECT	37.48 59.575 37.53 59.705 ;
		RECT	37.48 60.56 37.53 60.69 ;
		RECT	37.48 62.035 37.53 62.165 ;
		RECT	37.475 62.32 37.525 62.37 ;
		RECT	37.48 63.02 37.53 63.15 ;
		RECT	37.475 66.21 37.525 66.34 ;
		RECT	37.475 66.955 37.525 67.085 ;
		RECT	37.475 68.435 37.525 68.565 ;
		RECT	38.015 29.565 38.065 29.695 ;
		RECT	38.015 31.04 38.065 31.17 ;
		RECT	38.015 31.79 38.065 31.92 ;
		RECT	38.015 33.785 38.065 33.835 ;
		RECT	38.015 34.985 38.065 35.115 ;
		RECT	38.015 35.96 38.065 36.09 ;
		RECT	38.015 37.435 38.065 37.565 ;
		RECT	38.015 38.42 38.065 38.55 ;
		RECT	38.015 39.9 38.065 40.03 ;
		RECT	38.015 40.39 38.065 40.52 ;
		RECT	38.015 42.85 38.065 42.98 ;
		RECT	38.015 44.31 38.065 44.44 ;
		RECT	38.015 46.095 38.065 46.225 ;
		RECT	38.015 46.41 38.065 46.54 ;
		RECT	38.015 48.26 38.065 48.39 ;
		RECT	38.015 49.735 38.065 49.865 ;
		RECT	38.015 51.525 38.065 51.655 ;
		RECT	38.015 51.87 38.065 52 ;
		RECT	38.02 53.675 38.07 53.805 ;
		RECT	38.02 55.15 38.07 55.28 ;
		RECT	38.02 58.1 38.07 58.23 ;
		RECT	38.02 59.575 38.07 59.705 ;
		RECT	38.02 60.56 38.07 60.69 ;
		RECT	38.02 62.035 38.07 62.165 ;
		RECT	38.015 62.32 38.065 62.37 ;
		RECT	38.02 63.02 38.07 63.15 ;
		RECT	38.015 66.21 38.065 66.34 ;
		RECT	38.015 66.955 38.065 67.085 ;
		RECT	38.015 68.435 38.065 68.565 ;
		RECT	38.555 29.565 38.605 29.695 ;
		RECT	38.555 31.04 38.605 31.17 ;
		RECT	38.555 31.79 38.605 31.92 ;
		RECT	38.555 33.785 38.605 33.835 ;
		RECT	38.555 34.985 38.605 35.115 ;
		RECT	38.555 35.96 38.605 36.09 ;
		RECT	38.555 37.435 38.605 37.565 ;
		RECT	38.555 38.42 38.605 38.55 ;
		RECT	38.555 39.9 38.605 40.03 ;
		RECT	38.555 40.39 38.605 40.52 ;
		RECT	38.555 42.85 38.605 42.98 ;
		RECT	38.555 44.31 38.605 44.44 ;
		RECT	38.555 46.095 38.605 46.225 ;
		RECT	38.555 46.41 38.605 46.54 ;
		RECT	38.555 48.26 38.605 48.39 ;
		RECT	38.555 49.735 38.605 49.865 ;
		RECT	38.555 51.525 38.605 51.655 ;
		RECT	38.555 51.87 38.605 52 ;
		RECT	38.56 53.675 38.61 53.805 ;
		RECT	38.56 55.15 38.61 55.28 ;
		RECT	38.56 58.1 38.61 58.23 ;
		RECT	38.56 59.575 38.61 59.705 ;
		RECT	38.56 60.56 38.61 60.69 ;
		RECT	38.56 62.035 38.61 62.165 ;
		RECT	38.555 62.32 38.605 62.37 ;
		RECT	38.56 63.02 38.61 63.15 ;
		RECT	38.555 66.21 38.605 66.34 ;
		RECT	38.555 66.955 38.605 67.085 ;
		RECT	38.555 68.435 38.605 68.565 ;
		RECT	39.095 29.565 39.145 29.695 ;
		RECT	39.095 31.04 39.145 31.17 ;
		RECT	39.095 31.79 39.145 31.92 ;
		RECT	39.095 33.785 39.145 33.835 ;
		RECT	39.095 34.985 39.145 35.115 ;
		RECT	39.095 35.96 39.145 36.09 ;
		RECT	39.095 37.435 39.145 37.565 ;
		RECT	39.095 38.42 39.145 38.55 ;
		RECT	39.095 39.9 39.145 40.03 ;
		RECT	39.095 40.39 39.145 40.52 ;
		RECT	39.095 42.85 39.145 42.98 ;
		RECT	39.095 44.31 39.145 44.44 ;
		RECT	39.095 46.095 39.145 46.225 ;
		RECT	39.095 46.41 39.145 46.54 ;
		RECT	39.095 48.26 39.145 48.39 ;
		RECT	39.095 49.735 39.145 49.865 ;
		RECT	39.095 51.525 39.145 51.655 ;
		RECT	39.095 51.87 39.145 52 ;
		RECT	39.1 53.675 39.15 53.805 ;
		RECT	39.1 55.15 39.15 55.28 ;
		RECT	39.1 58.1 39.15 58.23 ;
		RECT	39.1 59.575 39.15 59.705 ;
		RECT	39.1 60.56 39.15 60.69 ;
		RECT	39.1 62.035 39.15 62.165 ;
		RECT	39.095 62.32 39.145 62.37 ;
		RECT	39.1 63.02 39.15 63.15 ;
		RECT	39.095 66.21 39.145 66.34 ;
		RECT	39.095 66.955 39.145 67.085 ;
		RECT	39.095 68.435 39.145 68.565 ;
		RECT	39.635 29.565 39.685 29.695 ;
		RECT	39.635 31.04 39.685 31.17 ;
		RECT	39.635 31.79 39.685 31.92 ;
		RECT	39.635 33.785 39.685 33.835 ;
		RECT	39.635 34.985 39.685 35.115 ;
		RECT	39.635 35.96 39.685 36.09 ;
		RECT	39.635 37.435 39.685 37.565 ;
		RECT	39.635 38.42 39.685 38.55 ;
		RECT	39.635 39.9 39.685 40.03 ;
		RECT	39.635 40.39 39.685 40.52 ;
		RECT	39.635 42.85 39.685 42.98 ;
		RECT	39.635 44.31 39.685 44.44 ;
		RECT	39.635 46.095 39.685 46.225 ;
		RECT	39.635 46.41 39.685 46.54 ;
		RECT	39.635 48.26 39.685 48.39 ;
		RECT	39.635 49.735 39.685 49.865 ;
		RECT	39.635 51.525 39.685 51.655 ;
		RECT	39.635 51.87 39.685 52 ;
		RECT	39.64 53.675 39.69 53.805 ;
		RECT	39.64 55.15 39.69 55.28 ;
		RECT	39.64 58.1 39.69 58.23 ;
		RECT	39.64 59.575 39.69 59.705 ;
		RECT	39.64 60.56 39.69 60.69 ;
		RECT	39.64 62.035 39.69 62.165 ;
		RECT	39.635 62.32 39.685 62.37 ;
		RECT	39.64 63.02 39.69 63.15 ;
		RECT	39.635 66.21 39.685 66.34 ;
		RECT	39.635 66.955 39.685 67.085 ;
		RECT	39.635 68.435 39.685 68.565 ;
		RECT	40.175 29.565 40.225 29.695 ;
		RECT	40.175 31.04 40.225 31.17 ;
		RECT	40.175 31.79 40.225 31.92 ;
		RECT	40.175 33.785 40.225 33.835 ;
		RECT	40.175 34.985 40.225 35.115 ;
		RECT	40.175 35.96 40.225 36.09 ;
		RECT	40.175 37.435 40.225 37.565 ;
		RECT	40.175 38.42 40.225 38.55 ;
		RECT	40.175 39.9 40.225 40.03 ;
		RECT	40.175 40.39 40.225 40.52 ;
		RECT	40.175 42.85 40.225 42.98 ;
		RECT	40.175 44.31 40.225 44.44 ;
		RECT	40.175 46.095 40.225 46.225 ;
		RECT	40.175 46.41 40.225 46.54 ;
		RECT	40.175 48.26 40.225 48.39 ;
		RECT	40.175 49.735 40.225 49.865 ;
		RECT	40.175 51.525 40.225 51.655 ;
		RECT	40.175 51.87 40.225 52 ;
		RECT	40.18 53.675 40.23 53.805 ;
		RECT	40.18 55.15 40.23 55.28 ;
		RECT	40.18 58.1 40.23 58.23 ;
		RECT	40.18 59.575 40.23 59.705 ;
		RECT	40.18 60.56 40.23 60.69 ;
		RECT	40.18 62.035 40.23 62.165 ;
		RECT	40.175 62.32 40.225 62.37 ;
		RECT	40.18 63.02 40.23 63.15 ;
		RECT	40.175 66.21 40.225 66.34 ;
		RECT	40.175 66.955 40.225 67.085 ;
		RECT	40.175 68.435 40.225 68.565 ;
		RECT	40.715 29.565 40.765 29.695 ;
		RECT	40.715 31.04 40.765 31.17 ;
		RECT	40.715 31.79 40.765 31.92 ;
		RECT	40.715 33.785 40.765 33.835 ;
		RECT	40.715 34.985 40.765 35.115 ;
		RECT	40.715 35.96 40.765 36.09 ;
		RECT	40.715 37.435 40.765 37.565 ;
		RECT	40.715 38.42 40.765 38.55 ;
		RECT	40.715 39.9 40.765 40.03 ;
		RECT	40.715 40.39 40.765 40.52 ;
		RECT	40.715 42.85 40.765 42.98 ;
		RECT	40.715 44.31 40.765 44.44 ;
		RECT	40.715 46.095 40.765 46.225 ;
		RECT	40.715 46.41 40.765 46.54 ;
		RECT	40.715 48.26 40.765 48.39 ;
		RECT	40.715 49.735 40.765 49.865 ;
		RECT	40.715 51.525 40.765 51.655 ;
		RECT	40.715 51.87 40.765 52 ;
		RECT	40.72 53.675 40.77 53.805 ;
		RECT	40.72 55.15 40.77 55.28 ;
		RECT	40.72 58.1 40.77 58.23 ;
		RECT	40.72 59.575 40.77 59.705 ;
		RECT	40.72 60.56 40.77 60.69 ;
		RECT	40.72 62.035 40.77 62.165 ;
		RECT	40.715 62.32 40.765 62.37 ;
		RECT	40.72 63.02 40.77 63.15 ;
		RECT	40.715 66.21 40.765 66.34 ;
		RECT	40.715 66.955 40.765 67.085 ;
		RECT	40.715 68.435 40.765 68.565 ;
		RECT	41.255 29.565 41.305 29.695 ;
		RECT	41.255 31.04 41.305 31.17 ;
		RECT	41.255 31.79 41.305 31.92 ;
		RECT	41.255 33.785 41.305 33.835 ;
		RECT	41.255 34.985 41.305 35.115 ;
		RECT	41.255 35.96 41.305 36.09 ;
		RECT	41.255 37.435 41.305 37.565 ;
		RECT	41.255 38.42 41.305 38.55 ;
		RECT	41.255 39.9 41.305 40.03 ;
		RECT	41.255 40.39 41.305 40.52 ;
		RECT	41.255 42.85 41.305 42.98 ;
		RECT	41.255 44.31 41.305 44.44 ;
		RECT	41.255 46.095 41.305 46.225 ;
		RECT	41.255 46.41 41.305 46.54 ;
		RECT	41.255 48.26 41.305 48.39 ;
		RECT	41.255 49.735 41.305 49.865 ;
		RECT	41.255 51.525 41.305 51.655 ;
		RECT	41.255 51.87 41.305 52 ;
		RECT	41.26 53.675 41.31 53.805 ;
		RECT	41.26 55.15 41.31 55.28 ;
		RECT	41.26 58.1 41.31 58.23 ;
		RECT	41.26 59.575 41.31 59.705 ;
		RECT	41.26 60.56 41.31 60.69 ;
		RECT	41.26 62.035 41.31 62.165 ;
		RECT	41.255 62.32 41.305 62.37 ;
		RECT	41.26 63.02 41.31 63.15 ;
		RECT	41.255 66.21 41.305 66.34 ;
		RECT	41.255 66.955 41.305 67.085 ;
		RECT	41.255 68.435 41.305 68.565 ;
		RECT	41.795 29.565 41.845 29.695 ;
		RECT	41.795 31.04 41.845 31.17 ;
		RECT	41.795 31.79 41.845 31.92 ;
		RECT	41.795 33.785 41.845 33.835 ;
		RECT	41.795 34.985 41.845 35.115 ;
		RECT	41.795 35.96 41.845 36.09 ;
		RECT	41.795 37.435 41.845 37.565 ;
		RECT	41.795 38.42 41.845 38.55 ;
		RECT	41.795 39.9 41.845 40.03 ;
		RECT	41.795 40.39 41.845 40.52 ;
		RECT	41.795 42.85 41.845 42.98 ;
		RECT	41.795 44.31 41.845 44.44 ;
		RECT	41.795 46.095 41.845 46.225 ;
		RECT	41.795 46.41 41.845 46.54 ;
		RECT	41.795 48.26 41.845 48.39 ;
		RECT	41.795 49.735 41.845 49.865 ;
		RECT	41.795 51.525 41.845 51.655 ;
		RECT	41.795 51.87 41.845 52 ;
		RECT	41.8 53.675 41.85 53.805 ;
		RECT	41.8 55.15 41.85 55.28 ;
		RECT	41.8 58.1 41.85 58.23 ;
		RECT	41.8 59.575 41.85 59.705 ;
		RECT	41.8 60.56 41.85 60.69 ;
		RECT	41.8 62.035 41.85 62.165 ;
		RECT	41.795 62.32 41.845 62.37 ;
		RECT	41.8 63.02 41.85 63.15 ;
		RECT	41.795 66.21 41.845 66.34 ;
		RECT	41.795 66.955 41.845 67.085 ;
		RECT	41.795 68.435 41.845 68.565 ;
		RECT	42.335 29.565 42.385 29.695 ;
		RECT	42.335 31.04 42.385 31.17 ;
		RECT	42.335 31.79 42.385 31.92 ;
		RECT	42.335 33.785 42.385 33.835 ;
		RECT	42.335 34.985 42.385 35.115 ;
		RECT	42.335 35.96 42.385 36.09 ;
		RECT	42.335 37.435 42.385 37.565 ;
		RECT	42.335 38.42 42.385 38.55 ;
		RECT	42.335 39.9 42.385 40.03 ;
		RECT	42.335 40.39 42.385 40.52 ;
		RECT	42.335 42.85 42.385 42.98 ;
		RECT	42.335 44.31 42.385 44.44 ;
		RECT	42.335 46.095 42.385 46.225 ;
		RECT	42.335 46.41 42.385 46.54 ;
		RECT	42.335 48.26 42.385 48.39 ;
		RECT	42.335 49.735 42.385 49.865 ;
		RECT	42.335 51.525 42.385 51.655 ;
		RECT	42.335 51.87 42.385 52 ;
		RECT	42.34 53.675 42.39 53.805 ;
		RECT	42.34 55.15 42.39 55.28 ;
		RECT	42.34 58.1 42.39 58.23 ;
		RECT	42.34 59.575 42.39 59.705 ;
		RECT	42.34 60.56 42.39 60.69 ;
		RECT	42.34 62.035 42.39 62.165 ;
		RECT	42.335 62.32 42.385 62.37 ;
		RECT	42.34 63.02 42.39 63.15 ;
		RECT	42.335 66.21 42.385 66.34 ;
		RECT	42.335 66.955 42.385 67.085 ;
		RECT	42.335 68.435 42.385 68.565 ;
		RECT	42.875 29.565 42.925 29.695 ;
		RECT	42.875 31.04 42.925 31.17 ;
		RECT	42.875 31.79 42.925 31.92 ;
		RECT	42.875 33.785 42.925 33.835 ;
		RECT	42.875 34.985 42.925 35.115 ;
		RECT	42.875 35.96 42.925 36.09 ;
		RECT	42.875 37.435 42.925 37.565 ;
		RECT	42.875 38.42 42.925 38.55 ;
		RECT	42.875 39.9 42.925 40.03 ;
		RECT	42.875 40.39 42.925 40.52 ;
		RECT	42.875 42.85 42.925 42.98 ;
		RECT	42.875 44.31 42.925 44.44 ;
		RECT	42.875 46.095 42.925 46.225 ;
		RECT	42.875 46.41 42.925 46.54 ;
		RECT	42.875 48.26 42.925 48.39 ;
		RECT	42.875 49.735 42.925 49.865 ;
		RECT	42.875 51.525 42.925 51.655 ;
		RECT	42.875 51.87 42.925 52 ;
		RECT	42.88 53.675 42.93 53.805 ;
		RECT	42.88 55.15 42.93 55.28 ;
		RECT	42.88 58.1 42.93 58.23 ;
		RECT	42.88 59.575 42.93 59.705 ;
		RECT	42.88 60.56 42.93 60.69 ;
		RECT	42.88 62.035 42.93 62.165 ;
		RECT	42.875 62.32 42.925 62.37 ;
		RECT	42.88 63.02 42.93 63.15 ;
		RECT	42.875 66.21 42.925 66.34 ;
		RECT	42.875 66.955 42.925 67.085 ;
		RECT	42.875 68.435 42.925 68.565 ;
		RECT	43.415 29.565 43.465 29.695 ;
		RECT	43.415 31.04 43.465 31.17 ;
		RECT	43.415 31.79 43.465 31.92 ;
		RECT	43.415 33.785 43.465 33.835 ;
		RECT	43.415 34.985 43.465 35.115 ;
		RECT	43.415 35.96 43.465 36.09 ;
		RECT	43.415 37.435 43.465 37.565 ;
		RECT	43.415 38.42 43.465 38.55 ;
		RECT	43.415 39.9 43.465 40.03 ;
		RECT	43.415 40.39 43.465 40.52 ;
		RECT	43.415 42.85 43.465 42.98 ;
		RECT	43.415 44.31 43.465 44.44 ;
		RECT	43.415 46.095 43.465 46.225 ;
		RECT	43.415 46.41 43.465 46.54 ;
		RECT	43.415 48.26 43.465 48.39 ;
		RECT	43.415 49.735 43.465 49.865 ;
		RECT	43.415 51.525 43.465 51.655 ;
		RECT	43.415 51.87 43.465 52 ;
		RECT	43.42 53.675 43.47 53.805 ;
		RECT	43.42 55.15 43.47 55.28 ;
		RECT	43.42 58.1 43.47 58.23 ;
		RECT	43.42 59.575 43.47 59.705 ;
		RECT	43.42 60.56 43.47 60.69 ;
		RECT	43.42 62.035 43.47 62.165 ;
		RECT	43.415 62.32 43.465 62.37 ;
		RECT	43.42 63.02 43.47 63.15 ;
		RECT	43.415 66.21 43.465 66.34 ;
		RECT	43.415 66.955 43.465 67.085 ;
		RECT	43.415 68.435 43.465 68.565 ;
		RECT	43.955 29.565 44.005 29.695 ;
		RECT	43.955 31.04 44.005 31.17 ;
		RECT	43.955 31.79 44.005 31.92 ;
		RECT	43.955 33.785 44.005 33.835 ;
		RECT	43.955 34.985 44.005 35.115 ;
		RECT	43.955 35.96 44.005 36.09 ;
		RECT	43.955 37.435 44.005 37.565 ;
		RECT	43.955 38.42 44.005 38.55 ;
		RECT	43.955 39.9 44.005 40.03 ;
		RECT	43.955 40.39 44.005 40.52 ;
		RECT	43.955 42.85 44.005 42.98 ;
		RECT	43.955 44.31 44.005 44.44 ;
		RECT	43.955 46.095 44.005 46.225 ;
		RECT	43.955 46.41 44.005 46.54 ;
		RECT	43.955 48.26 44.005 48.39 ;
		RECT	43.955 49.735 44.005 49.865 ;
		RECT	43.955 51.525 44.005 51.655 ;
		RECT	43.955 51.87 44.005 52 ;
		RECT	43.96 53.675 44.01 53.805 ;
		RECT	43.96 55.15 44.01 55.28 ;
		RECT	43.96 58.1 44.01 58.23 ;
		RECT	43.96 59.575 44.01 59.705 ;
		RECT	43.96 60.56 44.01 60.69 ;
		RECT	43.96 62.035 44.01 62.165 ;
		RECT	43.955 62.32 44.005 62.37 ;
		RECT	43.96 63.02 44.01 63.15 ;
		RECT	43.955 66.21 44.005 66.34 ;
		RECT	43.955 66.955 44.005 67.085 ;
		RECT	43.955 68.435 44.005 68.565 ;
		RECT	44.495 29.565 44.545 29.695 ;
		RECT	44.495 31.04 44.545 31.17 ;
		RECT	44.495 31.79 44.545 31.92 ;
		RECT	44.495 33.785 44.545 33.835 ;
		RECT	44.495 34.985 44.545 35.115 ;
		RECT	44.495 35.96 44.545 36.09 ;
		RECT	44.495 37.435 44.545 37.565 ;
		RECT	44.495 38.42 44.545 38.55 ;
		RECT	44.495 39.9 44.545 40.03 ;
		RECT	44.495 40.39 44.545 40.52 ;
		RECT	44.495 42.85 44.545 42.98 ;
		RECT	44.495 44.31 44.545 44.44 ;
		RECT	44.495 46.095 44.545 46.225 ;
		RECT	44.495 46.41 44.545 46.54 ;
		RECT	44.495 48.26 44.545 48.39 ;
		RECT	44.495 49.735 44.545 49.865 ;
		RECT	44.495 51.525 44.545 51.655 ;
		RECT	44.495 51.87 44.545 52 ;
		RECT	44.5 53.675 44.55 53.805 ;
		RECT	44.5 55.15 44.55 55.28 ;
		RECT	44.5 58.1 44.55 58.23 ;
		RECT	44.5 59.575 44.55 59.705 ;
		RECT	44.5 60.56 44.55 60.69 ;
		RECT	44.5 62.035 44.55 62.165 ;
		RECT	44.495 62.32 44.545 62.37 ;
		RECT	44.5 63.02 44.55 63.15 ;
		RECT	44.495 66.21 44.545 66.34 ;
		RECT	44.495 66.955 44.545 67.085 ;
		RECT	44.495 68.435 44.545 68.565 ;
		RECT	45.035 29.565 45.085 29.695 ;
		RECT	45.035 31.04 45.085 31.17 ;
		RECT	45.035 31.79 45.085 31.92 ;
		RECT	45.035 33.785 45.085 33.835 ;
		RECT	45.035 34.985 45.085 35.115 ;
		RECT	45.035 35.96 45.085 36.09 ;
		RECT	45.035 37.435 45.085 37.565 ;
		RECT	45.035 38.42 45.085 38.55 ;
		RECT	45.035 39.9 45.085 40.03 ;
		RECT	45.035 40.39 45.085 40.52 ;
		RECT	45.035 42.85 45.085 42.98 ;
		RECT	45.035 44.31 45.085 44.44 ;
		RECT	45.035 46.095 45.085 46.225 ;
		RECT	45.035 46.41 45.085 46.54 ;
		RECT	45.035 48.26 45.085 48.39 ;
		RECT	45.035 49.735 45.085 49.865 ;
		RECT	45.035 51.525 45.085 51.655 ;
		RECT	45.035 51.87 45.085 52 ;
		RECT	45.04 53.675 45.09 53.805 ;
		RECT	45.04 55.15 45.09 55.28 ;
		RECT	45.04 58.1 45.09 58.23 ;
		RECT	45.04 59.575 45.09 59.705 ;
		RECT	45.04 60.56 45.09 60.69 ;
		RECT	45.04 62.035 45.09 62.165 ;
		RECT	45.035 62.32 45.085 62.37 ;
		RECT	45.04 63.02 45.09 63.15 ;
		RECT	45.035 66.21 45.085 66.34 ;
		RECT	45.035 66.955 45.085 67.085 ;
		RECT	45.035 68.435 45.085 68.565 ;
		RECT	45.575 29.565 45.625 29.695 ;
		RECT	45.575 31.04 45.625 31.17 ;
		RECT	45.575 31.79 45.625 31.92 ;
		RECT	45.575 33.785 45.625 33.835 ;
		RECT	45.575 34.985 45.625 35.115 ;
		RECT	45.575 35.96 45.625 36.09 ;
		RECT	45.575 37.435 45.625 37.565 ;
		RECT	45.575 38.42 45.625 38.55 ;
		RECT	45.575 39.9 45.625 40.03 ;
		RECT	45.575 40.39 45.625 40.52 ;
		RECT	45.575 42.85 45.625 42.98 ;
		RECT	45.575 44.31 45.625 44.44 ;
		RECT	45.575 46.095 45.625 46.225 ;
		RECT	45.575 46.41 45.625 46.54 ;
		RECT	45.575 48.26 45.625 48.39 ;
		RECT	45.575 49.735 45.625 49.865 ;
		RECT	45.575 51.525 45.625 51.655 ;
		RECT	45.575 51.87 45.625 52 ;
		RECT	45.58 53.675 45.63 53.805 ;
		RECT	45.58 55.15 45.63 55.28 ;
		RECT	45.58 58.1 45.63 58.23 ;
		RECT	45.58 59.575 45.63 59.705 ;
		RECT	45.58 60.56 45.63 60.69 ;
		RECT	45.58 62.035 45.63 62.165 ;
		RECT	45.575 62.32 45.625 62.37 ;
		RECT	45.58 63.02 45.63 63.15 ;
		RECT	45.575 66.21 45.625 66.34 ;
		RECT	45.575 66.955 45.625 67.085 ;
		RECT	45.575 68.435 45.625 68.565 ;
		RECT	46.115 29.565 46.165 29.695 ;
		RECT	46.115 31.04 46.165 31.17 ;
		RECT	46.115 31.79 46.165 31.92 ;
		RECT	46.115 33.785 46.165 33.835 ;
		RECT	46.115 34.985 46.165 35.115 ;
		RECT	46.115 35.96 46.165 36.09 ;
		RECT	46.115 37.435 46.165 37.565 ;
		RECT	46.115 38.42 46.165 38.55 ;
		RECT	46.115 39.9 46.165 40.03 ;
		RECT	46.115 40.39 46.165 40.52 ;
		RECT	46.115 42.85 46.165 42.98 ;
		RECT	46.115 44.31 46.165 44.44 ;
		RECT	46.115 46.095 46.165 46.225 ;
		RECT	46.115 46.41 46.165 46.54 ;
		RECT	46.115 48.26 46.165 48.39 ;
		RECT	46.115 49.735 46.165 49.865 ;
		RECT	46.115 51.525 46.165 51.655 ;
		RECT	46.115 51.87 46.165 52 ;
		RECT	46.12 53.675 46.17 53.805 ;
		RECT	46.12 55.15 46.17 55.28 ;
		RECT	46.12 58.1 46.17 58.23 ;
		RECT	46.12 59.575 46.17 59.705 ;
		RECT	46.12 60.56 46.17 60.69 ;
		RECT	46.12 62.035 46.17 62.165 ;
		RECT	46.115 62.32 46.165 62.37 ;
		RECT	46.12 63.02 46.17 63.15 ;
		RECT	46.115 66.21 46.165 66.34 ;
		RECT	46.115 66.955 46.165 67.085 ;
		RECT	46.115 68.435 46.165 68.565 ;
		RECT	46.655 29.565 46.705 29.695 ;
		RECT	46.655 31.04 46.705 31.17 ;
		RECT	46.655 31.79 46.705 31.92 ;
		RECT	46.655 33.785 46.705 33.835 ;
		RECT	46.655 34.985 46.705 35.115 ;
		RECT	46.655 35.96 46.705 36.09 ;
		RECT	46.655 37.435 46.705 37.565 ;
		RECT	46.655 38.42 46.705 38.55 ;
		RECT	46.655 39.9 46.705 40.03 ;
		RECT	46.655 40.39 46.705 40.52 ;
		RECT	46.655 42.85 46.705 42.98 ;
		RECT	46.655 44.31 46.705 44.44 ;
		RECT	46.655 46.095 46.705 46.225 ;
		RECT	46.655 46.41 46.705 46.54 ;
		RECT	46.655 48.26 46.705 48.39 ;
		RECT	46.655 49.735 46.705 49.865 ;
		RECT	46.655 51.525 46.705 51.655 ;
		RECT	46.655 51.87 46.705 52 ;
		RECT	46.66 53.675 46.71 53.805 ;
		RECT	46.66 55.15 46.71 55.28 ;
		RECT	46.66 58.1 46.71 58.23 ;
		RECT	46.66 59.575 46.71 59.705 ;
		RECT	46.66 60.56 46.71 60.69 ;
		RECT	46.66 62.035 46.71 62.165 ;
		RECT	46.655 62.32 46.705 62.37 ;
		RECT	46.66 63.02 46.71 63.15 ;
		RECT	46.655 66.21 46.705 66.34 ;
		RECT	46.655 66.955 46.705 67.085 ;
		RECT	46.655 68.435 46.705 68.565 ;
		RECT	47.195 29.565 47.245 29.695 ;
		RECT	47.195 31.04 47.245 31.17 ;
		RECT	47.195 31.79 47.245 31.92 ;
		RECT	47.195 33.785 47.245 33.835 ;
		RECT	47.195 34.985 47.245 35.115 ;
		RECT	47.195 35.96 47.245 36.09 ;
		RECT	47.195 37.435 47.245 37.565 ;
		RECT	47.195 38.42 47.245 38.55 ;
		RECT	47.195 39.9 47.245 40.03 ;
		RECT	47.195 40.39 47.245 40.52 ;
		RECT	47.195 42.85 47.245 42.98 ;
		RECT	47.195 44.31 47.245 44.44 ;
		RECT	47.195 46.095 47.245 46.225 ;
		RECT	47.195 46.41 47.245 46.54 ;
		RECT	47.195 48.26 47.245 48.39 ;
		RECT	47.195 49.735 47.245 49.865 ;
		RECT	47.195 51.525 47.245 51.655 ;
		RECT	47.195 51.87 47.245 52 ;
		RECT	47.2 53.675 47.25 53.805 ;
		RECT	47.2 55.15 47.25 55.28 ;
		RECT	47.2 58.1 47.25 58.23 ;
		RECT	47.2 59.575 47.25 59.705 ;
		RECT	47.2 60.56 47.25 60.69 ;
		RECT	47.2 62.035 47.25 62.165 ;
		RECT	47.195 62.32 47.245 62.37 ;
		RECT	47.2 63.02 47.25 63.15 ;
		RECT	47.195 66.21 47.245 66.34 ;
		RECT	47.195 66.955 47.245 67.085 ;
		RECT	47.195 68.435 47.245 68.565 ;
		RECT	47.735 29.565 47.785 29.695 ;
		RECT	47.735 31.04 47.785 31.17 ;
		RECT	47.735 31.79 47.785 31.92 ;
		RECT	47.735 33.785 47.785 33.835 ;
		RECT	47.735 34.985 47.785 35.115 ;
		RECT	47.735 35.96 47.785 36.09 ;
		RECT	47.735 37.435 47.785 37.565 ;
		RECT	47.735 38.42 47.785 38.55 ;
		RECT	47.735 39.9 47.785 40.03 ;
		RECT	47.735 40.39 47.785 40.52 ;
		RECT	47.735 42.85 47.785 42.98 ;
		RECT	47.735 44.31 47.785 44.44 ;
		RECT	47.735 46.095 47.785 46.225 ;
		RECT	47.735 46.41 47.785 46.54 ;
		RECT	47.735 48.26 47.785 48.39 ;
		RECT	47.735 49.735 47.785 49.865 ;
		RECT	47.735 51.525 47.785 51.655 ;
		RECT	47.735 51.87 47.785 52 ;
		RECT	47.74 53.675 47.79 53.805 ;
		RECT	47.74 55.15 47.79 55.28 ;
		RECT	47.74 58.1 47.79 58.23 ;
		RECT	47.74 59.575 47.79 59.705 ;
		RECT	47.74 60.56 47.79 60.69 ;
		RECT	47.74 62.035 47.79 62.165 ;
		RECT	47.735 62.32 47.785 62.37 ;
		RECT	47.74 63.02 47.79 63.15 ;
		RECT	47.735 66.21 47.785 66.34 ;
		RECT	47.735 66.955 47.785 67.085 ;
		RECT	47.735 68.435 47.785 68.565 ;
		RECT	48.275 29.565 48.325 29.695 ;
		RECT	48.275 31.04 48.325 31.17 ;
		RECT	48.275 31.79 48.325 31.92 ;
		RECT	48.275 33.785 48.325 33.835 ;
		RECT	48.275 34.985 48.325 35.115 ;
		RECT	48.275 35.96 48.325 36.09 ;
		RECT	48.275 37.435 48.325 37.565 ;
		RECT	48.275 38.42 48.325 38.55 ;
		RECT	48.275 39.9 48.325 40.03 ;
		RECT	48.275 40.39 48.325 40.52 ;
		RECT	48.275 42.85 48.325 42.98 ;
		RECT	48.275 44.31 48.325 44.44 ;
		RECT	48.275 46.095 48.325 46.225 ;
		RECT	48.275 46.41 48.325 46.54 ;
		RECT	48.275 48.26 48.325 48.39 ;
		RECT	48.275 49.735 48.325 49.865 ;
		RECT	48.275 51.525 48.325 51.655 ;
		RECT	48.275 51.87 48.325 52 ;
		RECT	48.28 53.675 48.33 53.805 ;
		RECT	48.28 55.15 48.33 55.28 ;
		RECT	48.28 58.1 48.33 58.23 ;
		RECT	48.28 59.575 48.33 59.705 ;
		RECT	48.28 60.56 48.33 60.69 ;
		RECT	48.28 62.035 48.33 62.165 ;
		RECT	48.275 62.32 48.325 62.37 ;
		RECT	48.28 63.02 48.33 63.15 ;
		RECT	48.275 66.21 48.325 66.34 ;
		RECT	48.275 66.955 48.325 67.085 ;
		RECT	48.275 68.435 48.325 68.565 ;
		RECT	48.815 29.565 48.865 29.695 ;
		RECT	48.815 31.04 48.865 31.17 ;
		RECT	48.815 31.79 48.865 31.92 ;
		RECT	48.815 33.785 48.865 33.835 ;
		RECT	48.815 34.985 48.865 35.115 ;
		RECT	48.815 35.96 48.865 36.09 ;
		RECT	48.815 37.435 48.865 37.565 ;
		RECT	48.815 38.42 48.865 38.55 ;
		RECT	48.815 39.9 48.865 40.03 ;
		RECT	48.815 40.39 48.865 40.52 ;
		RECT	48.815 42.85 48.865 42.98 ;
		RECT	48.815 44.31 48.865 44.44 ;
		RECT	48.815 46.095 48.865 46.225 ;
		RECT	48.815 46.41 48.865 46.54 ;
		RECT	48.815 48.26 48.865 48.39 ;
		RECT	48.815 49.735 48.865 49.865 ;
		RECT	48.815 51.525 48.865 51.655 ;
		RECT	48.815 51.87 48.865 52 ;
		RECT	48.82 53.675 48.87 53.805 ;
		RECT	48.82 55.15 48.87 55.28 ;
		RECT	48.82 58.1 48.87 58.23 ;
		RECT	48.82 59.575 48.87 59.705 ;
		RECT	48.82 60.56 48.87 60.69 ;
		RECT	48.82 62.035 48.87 62.165 ;
		RECT	48.815 62.32 48.865 62.37 ;
		RECT	48.82 63.02 48.87 63.15 ;
		RECT	48.815 66.21 48.865 66.34 ;
		RECT	48.815 66.955 48.865 67.085 ;
		RECT	48.815 68.435 48.865 68.565 ;
		RECT	49.355 29.565 49.405 29.695 ;
		RECT	49.355 31.04 49.405 31.17 ;
		RECT	49.355 31.79 49.405 31.92 ;
		RECT	49.355 33.785 49.405 33.835 ;
		RECT	49.355 34.985 49.405 35.115 ;
		RECT	49.355 35.96 49.405 36.09 ;
		RECT	49.355 37.435 49.405 37.565 ;
		RECT	49.355 38.42 49.405 38.55 ;
		RECT	49.355 39.9 49.405 40.03 ;
		RECT	49.355 40.39 49.405 40.52 ;
		RECT	49.355 42.85 49.405 42.98 ;
		RECT	49.355 44.31 49.405 44.44 ;
		RECT	49.355 46.095 49.405 46.225 ;
		RECT	49.355 46.41 49.405 46.54 ;
		RECT	49.355 48.26 49.405 48.39 ;
		RECT	49.355 49.735 49.405 49.865 ;
		RECT	49.355 51.525 49.405 51.655 ;
		RECT	49.355 51.87 49.405 52 ;
		RECT	49.36 53.675 49.41 53.805 ;
		RECT	49.36 55.15 49.41 55.28 ;
		RECT	49.36 58.1 49.41 58.23 ;
		RECT	49.36 59.575 49.41 59.705 ;
		RECT	49.36 60.56 49.41 60.69 ;
		RECT	49.36 62.035 49.41 62.165 ;
		RECT	49.355 62.32 49.405 62.37 ;
		RECT	49.36 63.02 49.41 63.15 ;
		RECT	49.355 66.21 49.405 66.34 ;
		RECT	49.355 66.955 49.405 67.085 ;
		RECT	49.355 68.435 49.405 68.565 ;
		RECT	49.705 29.54 49.835 29.72 ;
		RECT	50.09 30.34 50.22 30.39 ;
		RECT	49.705 30.585 49.835 30.635 ;
		RECT	50.09 31.32 50.22 31.37 ;
		RECT	49.705 32.49 49.835 32.67 ;
		RECT	50.125 33.01 50.175 33.14 ;
		RECT	49.705 33.54 49.835 33.59 ;
		RECT	49.705 33.785 49.835 33.835 ;
		RECT	50.125 33.99 50.175 34.12 ;
		RECT	49.94 34.485 49.99 34.615 ;
		RECT	49.705 36.43 49.835 36.61 ;
		RECT	50.125 36.945 50.175 37.075 ;
		RECT	49.705 37.41 49.835 37.59 ;
		RECT	49.705 38.395 49.835 38.575 ;
		RECT	49.705 40.365 49.835 40.545 ;
		RECT	50.125 40.88 50.175 41.01 ;
		RECT	49.705 41.345 49.835 41.525 ;
		RECT	50.125 41.865 50.175 41.995 ;
		RECT	49.705 42.33 49.835 42.51 ;
		RECT	49.705 44.305 49.835 44.485 ;
		RECT	50.125 44.815 50.175 44.945 ;
		RECT	49.705 45.285 49.835 45.465 ;
		RECT	50.09 47.07 50.22 47.12 ;
		RECT	50.09 47.565 50.22 47.615 ;
		RECT	49.705 48.235 49.835 48.415 ;
		RECT	50.125 48.75 50.175 48.88 ;
		RECT	50.125 49.245 50.175 49.375 ;
		RECT	49.705 49.71 49.835 49.89 ;
		RECT	50.09 50.515 50.22 50.565 ;
		RECT	50.09 51.005 50.22 51.055 ;
		RECT	49.705 52.66 49.835 52.84 ;
		RECT	50.125 53.18 50.175 53.31 ;
		RECT	49.705 53.65 49.835 53.83 ;
		RECT	49.705 55.615 49.835 55.795 ;
		RECT	50.125 56.135 50.175 56.265 ;
		RECT	49.705 56.6 49.835 56.78 ;
		RECT	50.125 57.115 50.175 57.245 ;
		RECT	49.705 57.585 49.835 57.765 ;
		RECT	49.705 59.55 49.835 59.73 ;
		RECT	49.705 60.535 49.835 60.715 ;
		RECT	50.125 61.055 50.175 61.185 ;
		RECT	49.705 61.52 49.835 61.7 ;
		RECT	49.705 62.32 49.835 62.37 ;
		RECT	49.94 63.515 49.99 63.645 ;
		RECT	50.125 64.005 50.175 64.135 ;
		RECT	49.705 64.47 49.835 64.65 ;
		RECT	50.125 64.955 50.175 65.085 ;
		RECT	49.705 65.455 49.835 65.635 ;
		RECT	50.09 66.755 50.22 66.805 ;
		RECT	49.705 67.49 49.835 67.54 ;
		RECT	50.125 67.735 50.175 67.785 ;
		RECT	49.705 68.475 49.835 68.525 ;
	END

END rf2_256x19_wm0

END LIBRARY

