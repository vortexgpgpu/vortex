
module VX_front_end (
	input clk,    // Clock
	input reset,
	input icache_response_t icache_response,


	output icache_request_t icache_request,
	
);





endmodule