`include "VX_rop_define.vh"

module VX_rop_ds #(
    parameter CLUSTER_ID = 0,
    parameter NUM_LANES  = 4
) (
    input wire clk,
    input wire reset
    // TODO
);

    // TODO

endmodule