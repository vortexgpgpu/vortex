`ifndef VX_TEX_DEFINE_VH
`define VX_TEX_DEFINE_VH

`include "VX_define.vh"
`include "VX_tex_types.vh"

`IGNORE_WARNINGS_BEGIN
import VX_tex_types::*;
`IGNORE_WARNINGS_END

`endif
