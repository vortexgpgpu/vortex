`include "VX_raster_define.vh"

module VX_raster_unit #(  
    parameter CORE_ID = 0
) (
    input wire  clk,
    input wire  reset

    // TODO
);

    // TODO

endmodule