`ifndef VX_ROP_DEFINE_VH
`define VX_ROP_DEFINE_VH

`include "VX_define.vh"
`include "VX_rop_types.vh"

`IGNORE_WARNINGS_BEGIN
import VX_rop_types::*;
`IGNORE_WARNINGS_END

`endif
