`include "VX_rop_define.vh"

module VX_rop_logic #(
    // TODO
) (
    input wire clk,
    input wire reset
    // TODO
);

    // TODO

endmodule