`include "VX_rop_define.vh"

module VX_rop_ds #(
    parameter `STRING_TYPE INSTANCE_ID = "",
    parameter NUM_LANES = 4,
    parameter TAG_WIDTH = 1
) (
    input wire clk,
    input wire reset,
    
    // DCRs
    input rop_dcrs_t dcrs,

    // Handshake
    input wire                  valid_in,
    input wire [TAG_WIDTH-1:0]  tag_in,
    output wire                 ready_in,   
     
    output wire                 valid_out,
    output wire [TAG_WIDTH-1:0] tag_out,
    input wire                  ready_out,

    // Input values
    input wire [NUM_LANES-1:0]                          face,
    input wire [NUM_LANES-1:0][`ROP_DEPTH_BITS-1:0]     depth_ref,
    input wire [NUM_LANES-1:0][`ROP_DEPTH_BITS-1:0]     depth_val,
    input wire [NUM_LANES-1:0][`ROP_STENCIL_BITS-1:0]   stencil_val,    

    // Output values
    output wire [NUM_LANES-1:0][`ROP_DEPTH_BITS-1:0]    depth_out,        
    output wire [NUM_LANES-1:0][`ROP_STENCIL_BITS-1:0]  stencil_out,
    output wire [NUM_LANES-1:0]                         pass_out
); 
    `UNUSED_VAR (dcrs)

    wire stall = ~ready_out && valid_out;
    
    assign ready_in = ~stall;
    
    // Depth Test /////////////////////////////////////////////////////////////

    wire [NUM_LANES-1:0] dpass;

    for (genvar i = 0; i < NUM_LANES; ++i) begin
        VX_rop_compare #(
            .DATAW (`ROP_DEPTH_BITS)
        ) rop_compare_depth (
            .func   (dcrs.depth_func),
            .a      (depth_ref[i]),
            .b      (depth_val[i]),
            .result (dpass[i])
        );
    end

    // Stencil Test ///////////////////////////////////////////////////////////

    wire [NUM_LANES-1:0] spass;

    for (genvar i = 0; i < NUM_LANES; ++i) begin
        VX_rop_compare #(
            .DATAW (`ROP_STENCIL_BITS)
        ) rop_compare_stencil (
            .func   (dcrs.stencil_func[face[i]]),
            .a      (dcrs.stencil_ref[face[i]] & dcrs.stencil_mask[face[i]]),
            .b      (stencil_val[i] & dcrs.stencil_mask[face[i]]),
            .result (spass[i])
        );
    end  

    ///////////////////////////////////////////////////////////////////////////

    wire valid_in_s;
    wire [NUM_LANES-1:0] face_s;
    wire [NUM_LANES-1:0] dpass_s, spass_s;
    wire [NUM_LANES-1:0][`ROP_DEPTH_BITS-1:0] depth_ref_s, depth_val_s;
    wire [NUM_LANES-1:0][`ROP_STENCIL_BITS-1:0] stencil_val_s;
    wire [TAG_WIDTH-1:0] tag_in_s;
    
    VX_pipe_register #(
        .DATAW	(1 + NUM_LANES * (1 + 1 + 1 + 2 * `ROP_DEPTH_BITS + `ROP_STENCIL_BITS) + TAG_WIDTH),
        .RESETW (1),
        .DEPTH  (2)
    ) pipe_reg1 (
        .clk      (clk),
        .reset    (reset),
        .enable   (~stall),
        .data_in  ({valid_in,   face,   dpass,   spass,   depth_ref,   depth_val,   stencil_val,   tag_in}),
        .data_out ({valid_in_s, face_s, dpass_s, spass_s, depth_ref_s, depth_val_s, stencil_val_s, tag_in_s})
    );

    // Stencil Operation //////////////////////////////////////////////////////

    wire [NUM_LANES-1:0][`ROP_STENCIL_BITS-1:0] stencil_result;

    for (genvar i = 0; i < NUM_LANES; ++i) begin
        wire [`ROP_STENCIL_OP_BITS-1:0] stencil_op;
        assign stencil_op = spass_s[i] ? (dpass_s[i] ? dcrs.stencil_zpass[face_s[i]]
                                                     : dcrs.stencil_zfail[face_s[i]])
                                       : dcrs.stencil_fail[face_s[i]];
        VX_rop_stencil_op #(
            .DATAW (`ROP_STENCIL_BITS)
        ) rop_stencil_op (
            .stencil_op     (stencil_op),
            .stencil_ref    (dcrs.stencil_ref[face_s[i]]),
            .stencil_val    (stencil_val_s[i]),
            .stencil_result (stencil_result[i])
        );
    end

    ///////////////////////////////////////////////////////////////////////////

    wire [NUM_LANES-1:0][`ROP_DEPTH_BITS-1:0]   depth_write;
    wire [NUM_LANES-1:0][`ROP_STENCIL_BITS-1:0] stencil_write;
    wire [NUM_LANES-1:0] pass;

    for (genvar i = 0; i < NUM_LANES; ++i) begin
        assign depth_write[i] = (dpass_s[i] && dcrs.depth_writemask) ? depth_ref_s[i] : depth_val_s[i];
        for (genvar j = 0; j < `ROP_STENCIL_BITS; ++j) begin
            assign stencil_write[i][j] = dcrs.stencil_writemask[face_s[i]][j] ? stencil_result[i][j] : stencil_val_s[i][j];
        end
    end

    assign pass = spass_s & dpass_s;

    // Output /////////////////////////////////////////////////////////////////

    VX_pipe_register #(
        .DATAW	(1 + TAG_WIDTH + NUM_LANES * (`ROP_DEPTH_BITS + `ROP_STENCIL_BITS + 1)),
        .RESETW (1)
    ) pipe_reg2 (
        .clk      (clk),
        .reset    (reset),
        .enable   (~stall),
        .data_in  ({valid_in_s, tag_in_s, depth_write, stencil_write, pass}),
        .data_out ({valid_out,  tag_out,  depth_out,   stencil_out,   pass_out})
    );

endmodule
