`ifndef VX_CACHE_CONFIG
`define VX_CACHE_CONFIG

`include "../VX_define.vh"

//                                data         tid                   rd  wb    warp_num  read write
`define MRVQ_METADATA_SIZE      (`WORD_SIZE + `LOG2UP(NUM_REQUESTS) + 5 + 2 + (`NW_BITS) + 3 + 3)

//                               rd  wb   warp_num  read write + reqs
`define REQ_INST_META_SIZE      (5 + 2 + (`NW_BITS) + 3 + 3 + `LOG2UP(NUM_REQUESTS))

`define WORD_SIZE               (8 * WORD_SIZE_BYTES)
`define WORD_SIZE_RNG           (`WORD_SIZE)-1:0

// 128
`define BANK_SIZE_BYTES         (CACHE_SIZE_BYTES / NUM_BANKS)      

// 8
`define BANK_LINE_COUNT         (`BANK_SIZE_BYTES / BANK_LINE_SIZE_BYTES)
// 4
`define BANK_LINE_WORDS         (BANK_LINE_SIZE_BYTES / WORD_SIZE_BYTES)

// Offset is fixed
`define OFFSET_ADDR_BITS        2
`define OFFSET_SIZE_END         1
`define OFFSET_ADDR_START       0
`define OFFSET_ADDR_END         1
`define OFFSET_ADDR_RNG         `OFFSET_ADDR_END:`OFFSET_ADDR_START
`define OFFSET_SIZE_RNG         `OFFSET_SIZE_END:0

// 2
`define WORD_SELECT_BITS        (`LOG2UP(`BANK_LINE_WORDS))
// 2
`define WORD_SELECT_SIZE_END    (`WORD_SELECT_BITS)
// 2
`define WORD_SELECT_ADDR_START  (1+`OFFSET_ADDR_END)
// 3
`define WORD_SELECT_ADDR_END    (`WORD_SELECT_SIZE_END+`OFFSET_ADDR_END)
// 3:2
`define WORD_SELECT_ADDR_RNG    `WORD_SELECT_ADDR_END:`WORD_SELECT_ADDR_START

// 3
`define BANK_SELECT_BITS        (`LOG2UP(NUM_BANKS))
// 3
`define BANK_SELECT_SIZE_END    (`BANK_SELECT_BITS)
// 4
`define BANK_SELECT_ADDR_START  (1+`WORD_SELECT_ADDR_END)
// 6
`define BANK_SELECT_ADDR_END    (`BANK_SELECT_SIZE_END+`BANK_SELECT_ADDR_START-1)
// 6:4
`define BANK_SELECT_ADDR_RNG    `BANK_SELECT_ADDR_END:`BANK_SELECT_ADDR_START

// 3
`define LINE_SELECT_BITS        (`LOG2UP(`BANK_LINE_COUNT))
// 7
`define LINE_SELECT_ADDR_START  (1+`BANK_SELECT_ADDR_END)
// 9
`define LINE_SELECT_ADDR_END    (`LINE_SELECT_BITS+`LINE_SELECT_ADDR_START-1)
// 9:7
`define LINE_SELECT_ADDR_RNG    `LINE_SELECT_ADDR_END:`LINE_SELECT_ADDR_START

// 10
`define TAG_SELECT_ADDR_START   (1+`LINE_SELECT_ADDR_END)
// 31:10
`define TAG_SELECT_ADDR_RNG     31:`TAG_SELECT_ADDR_START
// 22
`define TAG_SELECT_BITS         (32-`TAG_SELECT_ADDR_START)

`define TAG_LINE_SELECT_BITS    (`TAG_SELECT_BITS+`LINE_SELECT_BITS)

`define BASE_ADDR_MASK          (~((1<<(`WORD_SELECT_ADDR_END+1))-1))

`endif
