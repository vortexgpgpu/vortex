`include "VX_define.vh"

module vortex_afu #(
	parameter AXI_DATA_WIDTH     = `VX_MEM_DATA_WIDTH,
    parameter AXI_ADDR_WIDTH     = `VX_MEM_ADDR_WIDTH,
    parameter AXI_TID_WIDTH      = 12,
    parameter AXI_STROBE_WIDTH   = `VX_MEM_BYTEEN_WIDTH,
	parameter AXI_DCR_ADDR_WIDTH = `VX_DCR_ADDR_WIDTH,
    parameter AXI_DCR_DATA_WIDTH = `VX_DCR_DATA_WIDTH    
) (
	// System signals
	input  wire  ap_clk,
	input  wire  ap_rst_n,
	
	// AXI4 master interface 
	output wire                                 m_axi_gmem_AWVALID,
	input  wire                                 m_axi_gmem_AWREADY,
	output wire [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m_axi_gmem_AWADDR,
	output wire [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m_axi_gmem_AWID,
	output wire [7:0]                           m_axi_gmem_AWLEN,
	output wire [2:0]                           m_axi_gmem_AWSIZE,
	// Tie-off AXI4 transaction options that are not being used.
	output wire [1:0]                           m_axi_gmem_AWBURST,
	output wire [1:0]                           m_axi_gmem_AWLOCK,
	output wire [3:0]                           m_axi_gmem_AWCACHE,
	output wire [2:0]                           m_axi_gmem_AWPROT,
	output wire [3:0]                           m_axi_gmem_AWQOS,
	output wire [3:0]                           m_axi_gmem_AWREGION,
	output wire                                 m_axi_gmem_WVALID,
	input  wire                                 m_axi_gmem_WREADY,
	output wire [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m_axi_gmem_WDATA,
	output wire [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m_axi_gmem_WSTRB,
	output wire                                 m_axi_gmem_WLAST,
	output wire                                 m_axi_gmem_ARVALID,
	input  wire                                 m_axi_gmem_ARREADY,
	output wire [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m_axi_gmem_ARADDR,
	output wire [C_M_AXI_GMEM_ID_WIDTH-1:0]     m_axi_gmem_ARID,
	output wire [7:0]                           m_axi_gmem_ARLEN,
	output wire [2:0]                           m_axi_gmem_ARSIZE,
	output wire [1:0]                           m_axi_gmem_ARBURST,
	output wire [1:0]                           m_axi_gmem_ARLOCK,
	output wire [3:0]                           m_axi_gmem_ARCACHE,
	output wire [2:0]                           m_axi_gmem_ARPROT,
	output wire [3:0]                           m_axi_gmem_ARQOS,
	output wire [3:0]                           m_axi_gmem_ARREGION,
	input  wire                                 m_axi_gmem_RVALID,
	output wire                                 m_axi_gmem_RREADY,
	input  wire [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m_axi_gmem_RDATA,
	input  wire                                 m_axi_gmem_RLAST,
	input  wire [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m_axi_gmem_RID,
	input  wire [1:0]                           m_axi_gmem_RRESP,
	input  wire                                 m_axi_gmem_BVALID,
	output wire                                 m_axi_gmem_BREADY,
	input  wire [1:0]                           m_axi_gmem_BRESP,
	input  wire [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m_axi_gmem_BID,

	// AXI4-Lite slave interface
	input  wire                                    s_axi_control_AWVALID,
	output wire                                    s_axi_control_AWREADY,
	input  wire [C_S_AXI_CONTROL_ADDR_WIDTH-1:0]   s_axi_control_AWADDR,
	input  wire                                    s_axi_control_WVALID,
	output wire                                    s_axi_control_WREADY,
	input  wire [C_S_AXI_CONTROL_DATA_WIDTH-1:0]   s_axi_control_WDATA,
	input  wire [C_S_AXI_CONTROL_DATA_WIDTH/8-1:0] s_axi_control_WSTRB,
	input  wire                                    s_axi_control_ARVALID,
	output wire                                    s_axi_control_ARREADY,
	input  wire [C_S_AXI_CONTROL_ADDR_WIDTH-1:0]   s_axi_control_ARADDR,
	output wire                                    s_axi_control_RVALID,
	input  wire                                    s_axi_control_RREADY,
	output wire [C_S_AXI_CONTROL_DATA_WIDTH-1:0]   s_axi_control_RDATA,
	output wire [1:0]                              s_axi_control_RRESP,
	output wire                                    s_axi_control_BVALID,
	input  wire                                    s_axi_control_BREADY,
	output wire [1:0]                              s_axi_control_BRESP
);

	Vortex_axi #(
		.AXI_DATA_WIDTH     (AXI_DATA_WIDTH),
		.AXI_ADDR_WIDTH     (AXI_ADDR_WIDTH),
		.AXI_TID_WIDTH      (AXI_TID_WIDTH),
		.AXI_STROBE_WIDTH   (AXI_STROBE_WIDTH),
		.AXI_DCR_ADDR_WIDTH (AXI_DCR_ADDR_WIDTH),
		.AXI_DCR_DATA_WIDTH (AXI_DCR_DATA_WIDTH)
	) inst (
		.clk(clk),
		.reset(reset),
		.m_axi_awid(m_axi_awid),
		.m_axi_awaddr(m_axi_awaddr),
		.m_axi_awlen(m_axi_awlen),
		.m_axi_awsize(m_axi_awsize),
		.m_axi_awburst(m_axi_awburst),
		.m_axi_awlock(m_axi_awlock),
		.m_axi_awcache(m_axi_awcache),
		.m_axi_awprot(m_axi_awprot),
		.m_axi_awqos(m_axi_awqos),
		.m_axi_awvalid(m_axi_awvalid),
		.m_axi_awready(m_axi_awready),
		.m_axi_wdata(m_axi_wdata),
		.m_axi_wstrb(m_axi_wstrb),
		.m_axi_wlast(m_axi_wlast),
		.m_axi_wvalid(m_axi_wvalid),
		.m_axi_wready(m_axi_wready),
		.m_axi_bid(m_axi_bid),
		.m_axi_bresp(m_axi_bresp),
		.m_axi_bvalid(m_axi_bvalid),
		.m_axi_bready(m_axi_bready),
		.m_axi_arid(m_axi_arid),
		.m_axi_araddr(m_axi_araddr),
		.m_axi_arlen(m_axi_arlen),
		.m_axi_arsize(m_axi_arsize),
		.m_axi_arburst(m_axi_arburst),
		.m_axi_arlock(m_axi_arlock),
		.m_axi_arcache(m_axi_arcache),
		.m_axi_arprot(m_axi_arprot),
		.m_axi_arqos(m_axi_arqos),
		.m_axi_arvalid(m_axi_arvalid),
		.m_axi_arready(m_axi_arready),
		.m_axi_rid(m_axi_rid),
		.m_axi_rdata(m_axi_rdata),
		.m_axi_rresp(m_axi_rresp),
		.m_axi_rlast(m_axi_rlast),
		.m_axi_rvalid(m_axi_rvalid),
		.m_axi_rready(m_axi_rready),
		.busy(busy)
	);
	
endmodule