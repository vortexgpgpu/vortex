`include "VX_raster_define.vh"

module VX_raster_fetch #( 
    // TODO
) (
    input wire clk,
    input wire reset
    // TODO
);

    // TODO

endmodule