`include "VX_rop_define.vh"

import VX_rop_types::*;

module VX_rop_req_switch #(
    // TODO
) (
    input wire clk,
    input wire reset
    // TODO
);

    // TODO

endmodule
