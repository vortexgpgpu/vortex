`ifndef __VORTEX_AFU__
`define __VORTEX_AFU__

`include "ccip_if_pkg.sv"

`define PLATFORM_PROVIDES_LOCAL_MEMORY
`define PLATFORM_PARAM_LOCAL_MEMORY_ADDR_WIDTH      27
`define PLATFORM_PARAM_LOCAL_MEMORY_DATA_WIDTH      512
`define PLATFORM_PARAM_LOCAL_MEMORY_BURST_CNT_WIDTH 4

`include "local_mem_cfg_pkg.sv"

`define AFU_ACCEL_NAME "vortex_afu"
`define AFU_ACCEL_UUID 128'h35f9452b_25c2_434c_93d5_6f8c60db361c
`define AFU_IMAGE_CMD_TYPE_CLFLUSH 4
`define AFU_IMAGE_CMD_TYPE_READ 1
`define AFU_IMAGE_CMD_TYPE_RUN 3
`define AFU_IMAGE_CMD_TYPE_WRITE 2
`define AFU_IMAGE_MMIO_CSR_CMD 10
`define AFU_IMAGE_MMIO_CSR_DATA_SIZE 12
`define AFU_IMAGE_MMIO_CSR_IO_ADDR 14
`define AFU_IMAGE_MMIO_CSR_MEM_ADDR 16
`define AFU_IMAGE_MMIO_CSR_STATUS 18
`define AFU_IMAGE_MMIO_CSR_SCOPE_CMD  20
`define AFU_IMAGE_MMIO_CSR_SCOPE_DATA 22
`define AFU_IMAGE_POWER 0
`define AFU_TOP_IFC "ccip_std_afu_avalon_mm"

`endif