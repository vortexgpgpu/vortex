`include "VX_raster_define.vh"

module VX_raster_slice #(  
    // TODO
) (
    input wire clk,
    input wire reset
    // TODO
);

    // TODO

endmodule