`include "VX_define.vh"

module VX_instr_sched #(
    parameter CORE_ID = 0
) (
    input wire clk,
    input wire reset,

    // inputs
    VX_decode_if  decode_if,  

    // outputs
    VX_instr_sched_if  instr_sched_if
);

    `UNUSED_PARAM (CORE_ID)
    
    localparam DATAW   = `NUM_THREADS + 32 + `EX_BITS + `OP_BITS + `FRM_BITS + 1 + (`NR_BITS * 4) + 32 + 1 + 1 + `NUM_REGS;
    localparam SIZE    = 3;
    localparam ADDRW   = $clog2(SIZE);
    localparam NWARPSW = $clog2(`NUM_WARPS+1);

    reg [`NUM_WARPS-1:0][ADDRW-1:0] used_r;
    reg [`NUM_WARPS-1:0] full_r, empty_r, alm_empty_r;
    
    wire [`NUM_WARPS-1:0] q_full, q_empty, q_alm_empty;
    wire [DATAW-1:0] q_data_in;
    wire [`NUM_WARPS-1:0][DATAW-1:0] q_data_prev;    
    reg [`NUM_WARPS-1:0][DATAW-1:0] q_data_out;

    wire enq_fire = decode_if.valid && decode_if.ready;
    wire deq_fire = instr_sched_if.valid && instr_sched_if.ready;

    for (genvar i = 0; i < `NUM_WARPS; ++i) begin

        wire writing = enq_fire && (i == decode_if.wid); 
        wire reading = deq_fire && (i == instr_sched_if.wid);

        wire is_head_ptr = empty_r[i] || (alm_empty_r[i] && reading);

        VX_skid_buffer #(
            .DATAW (DATAW)
        ) queue (
            .clk      (clk),
            .reset    (reset),
            .valid_in (writing && !is_head_ptr),
            .data_in  (q_data_in),            
            .ready_out(reading),
            .data_out (q_data_prev[i]),            
            `UNUSED_PIN (ready_in),
            `UNUSED_PIN (valid_out)
        );

        always @(posedge clk) begin
            if (reset) begin            
                used_r[i]      <= 0;
                full_r[i]      <= 0; 
                empty_r[i]     <= 1; 
                alm_empty_r[i] <= 1;
            end else begin  
                if (writing) begin
                    if (!reading) begin
                        empty_r[i] <= 0;
                        if (used_r[i] == 1)
                            alm_empty_r[i] <= 0;
                        if (used_r[i] == ADDRW'(SIZE-1))
                            full_r[i] <= 1;
                    end
                end else if (reading) begin
                    full_r[i] <= 0; 
                    if (used_r[i] == ADDRW'(1))
                        empty_r[i] <= 1;
                    if (used_r[i] == ADDRW'(2))
                        alm_empty_r[i] <= 1;
                end
                used_r[i] <= used_r[i] + ADDRW'($signed(2'(writing) - 2'(reading)));
            end 

            if (writing && is_head_ptr) begin                                                       
                q_data_out[i] <= q_data_in;
            end else if (reading) begin
                q_data_out[i] <= q_data_prev[i];
            end                  
        end
        
        assign q_full[i]      = full_r[i];
        assign q_empty[i]     = empty_r[i];
        assign q_alm_empty[i] = alm_empty_r[i];
    end

    ///////////////////////////////////////////////////////////////////////////

    reg [`NUM_WARPS-1:0] valid_table, valid_table_n;
    reg [`NUM_WARPS-1:0] schedule_table, schedule_table_n;
    reg [`NW_BITS-1:0] deq_wid, deq_wid_n;
    reg deq_valid, deq_valid_n;
    reg [DATAW-1:0] deq_instr, deq_instr_n;
    reg [NWARPSW-1:0] num_warps;

    // calculate valid table
    always @(*) begin
        valid_table_n = valid_table;        
        if (deq_fire) begin
            valid_table_n[deq_wid] = !q_alm_empty[deq_wid];
        end
        if (enq_fire) begin
            valid_table_n[decode_if.wid] = 1;
        end
    end

    // schedule the next instruction to issue
    always @(*) begin
        if (num_warps > 1) begin
            deq_valid_n = 1;
            deq_wid_n   = 'x;        
            deq_instr_n = 'x;
            for (integer i = `NUM_WARPS-1; i >= 0; --i) begin
                if (schedule_table[i]) begin
                    deq_wid_n   = `NW_BITS'(i);          
                    deq_instr_n = q_data_out[i];
                end
            end
        end else if (1 == num_warps && !(deq_fire && q_alm_empty[deq_wid])) begin
            deq_valid_n = 1;
            deq_wid_n   = deq_wid;
            deq_instr_n = deq_fire ? q_data_prev[deq_wid] : q_data_out[deq_wid];
        end else begin
            deq_valid_n = enq_fire;
            deq_wid_n   = decode_if.wid;
            deq_instr_n = q_data_in;  
        end   
    end

    // do round-robin scheduling with multiple active warps
    always @(*) begin
        if (1 == $countones(schedule_table) 
         || (num_warps < 2)) begin
            schedule_table_n = valid_table_n;            
        end else begin
            schedule_table_n = schedule_table;
        end
        schedule_table_n[deq_wid_n] = 0;
    end

    wire warp_added   = enq_fire && q_empty[decode_if.wid];
    wire warp_removed = deq_fire && ~(enq_fire && decode_if.wid == deq_wid) && q_alm_empty[deq_wid];
    
    always @(posedge clk) begin
        if (reset)  begin            
            valid_table    <= 0;
            deq_valid      <= 0;  
            num_warps      <= 0;         
        end else begin
            valid_table    <= valid_table_n;            
            deq_valid      <= deq_valid_n;
            schedule_table <= schedule_table_n;

            if (warp_added && !warp_removed) begin
                num_warps <= num_warps + NWARPSW'(1);
            end else if (warp_removed && !warp_added) begin
                num_warps <= num_warps - NWARPSW'(1);                
            end
        end
            
        deq_wid   <= deq_wid_n;
        deq_instr <= deq_instr_n;     
    end
    
    assign decode_if.ready = ~q_full[decode_if.wid];
    assign q_data_in = {decode_if.tmask, 
                        decode_if.PC, 
                        decode_if.ex_type, 
                        decode_if.op_type, 
                        decode_if.op_mod, 
                        decode_if.wb, 
                        decode_if.rd, 
                        decode_if.rs1, 
                        decode_if.rs2, 
                        decode_if.rs3, 
                        decode_if.imm, 
                        decode_if.use_PC, 
                        decode_if.use_imm,
                        decode_if.used_regs};

    assign instr_sched_if.valid = deq_valid;
    assign instr_sched_if.wid   = deq_wid;
    assign instr_sched_if.wid_n = deq_wid_n;
    assign {instr_sched_if.tmask, 
            instr_sched_if.PC, 
            instr_sched_if.ex_type, 
            instr_sched_if.op_type, 
            instr_sched_if.op_mod, 
            instr_sched_if.wb, 
            instr_sched_if.rd, 
            instr_sched_if.rs1, 
            instr_sched_if.rs2, 
            instr_sched_if.rs3, 
            instr_sched_if.imm, 
            instr_sched_if.use_PC, 
            instr_sched_if.use_imm, 
            instr_sched_if.used_regs} = deq_instr;

endmodule