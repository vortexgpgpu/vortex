`include "VX_rop_define.vh"

module VX_rop_blend #(  
    parameter CORE_ID = 0
    // TODO
) (
    input wire clk,
    input wire reset
    // TODO
);

    // TODO

endmodule