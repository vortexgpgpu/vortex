`timescale 1ns/1ps

module VX_tb_divide();

    `ifdef TRACE
    initial
    begin
    $dumpfile("trace.vcd");
    $dumpvars(0,test);
    end
    `endif

    reg clk;
    reg rst;

    reg [31:0] numer, denom;

    wire [31:0] o_div[0:7], o_rem[0:7];

    genvar i;
    generate
        for (i = 0; i < 8; i++) begin : div_loop
            VX_divide#(
                .WIDTHN(32),
                .WIDTHD(32),
                .PIPELINE(i)
            ) div(
                .clock(clk),
                .aclr(rst),
                .clken(1'b1),
                .numer(numer),
                .denom(denom),
                .quotient(o_div[i]),
                .remainder(o_rem[i])
            );
        end
    endgenerate

    initial begin
        clk = 0; rst = 0;

        numer = 56;
        denom = 11;

        $display("56 / 11 #0");
        if (o_div[0] != 5 || o_rem[0] != 1) begin
            $display("PIPE0: div=", o_div[0], " rem=", o_rem[0]);
            $display("expected 5,1 EXITING");
            $finish();
        end

        if (o_div[1] != 1'bx || o_rem[1] != 1'bx) begin
            $display("PIPE1: div=", o_div[1], " rem=", o_rem[1]);
            $display("expected x,x EXITING");
            $finish();
        end

        if (o_div[2] != 1'bx || o_rem[2] != 1'bx) begin
            $display("PIPE2: div=", o_div[2], " rem=", o_rem[2]);
            $display("expected x,x EXITING");
            $finish();
        end

        if (o_div[3] != 1'bx || o_rem[3] != 1'bx) begin
            $display("PIPE3: div=", o_div[3], " rem=", o_rem[3]);
            $display("expected x,x EXITING");
            $finish();
        end

        #2;

        $display("56 / 11 #2");
         if (o_div[0] != 5 || o_rem[0] != 1) begin
            $display("PIPE0: div=", o_div[0], " rem=", o_rem[0]);
            $display("expected 5,1, EXITING");
            $finish();
        end

        if (o_div[1] != 5 || o_rem[1] != 1) begin
            $display("PIPE1: div=", o_div[1], " rem=", o_rem[1]);
            $display("expected 5,1 EXITING");
            $finish();
        end

        if (o_div[2] != 1'bx || o_rem[2] != 1'bx) begin
            $display("PIPE2: div=", o_div[2], " rem=", o_rem[2]);
            $display("expected x,x EXITING");
            $finish();
        end

        if (o_div[3] != 1'bx || o_rem[3] != 1'bx) begin
            $display("PIPE3: div=", o_div[3], " rem=", o_rem[3]);
            $display("expected x,x EXITING");
            $finish();
        end

        #2;

        $display("56 / 11 #4");
        if (o_div[0] != 5 || o_rem[0] != 1) begin
            $display("PIPE0: div=", o_div[0], " rem=", o_rem[0]);
            $display("expected 5,1 EXITING");
            $finish();
        end

        if (o_div[1] != 5 || o_rem[1] != 1) begin
            $display("PIPE1: div=", o_div[1], " rem=", o_rem[1]);
            $display("expected 5,1 EXITING");
            $finish();
        end

        if (o_div[2] != 5 || o_rem[2] != 1) begin
            $display("PIPE2: div=", o_div[2], " rem=", o_rem[2]);
            $display("expected 5,1 EXITING");
            $finish();
        end

        if (o_div[3] != 1'bx || o_rem[3] != 1'bx) begin
            $display("PIPE3: div=", o_div[3], " rem=", o_rem[3]);
            $display("expected x,x EXITING");
            $finish();
        end

        #2;

        $display("56 / 11 #6");

        if (o_div[0] != 5 || o_rem[0] != 1) begin
            $display("PIPE0: div=", o_div[0], " rem=", o_rem[0]);
            $display("expected 5,1 EXITING");
            $finish();
        end

        if (o_div[1] != 5 || o_rem[1] != 1) begin
            $display("PIPE1: div=", o_div[1], " rem=", o_rem[1]);
            $display("expected 5,1 EXITING");
            $finish();
        end

        if (o_div[2] != 5 || o_rem[2] != 1) begin
            $display("PIPE2: div=", o_div[2], " rem=", o_rem[2]);
            $display("expected 5,1 EXITING");
            $finish();
        end

        if (o_div[3] != 5 || o_rem[3] != 1) begin
            $display("PIPE3: div=", o_div[3], " rem=", o_rem[3]);
            $display("expected 5,1 EXITING");
            $finish();
        end

        $display("PASS");

        $finish();
    end

    always #1
        clk = ~clk;

endmodule: VX_tb_divide