`include "VX_raster_define.vh"

module VX_raster_req_switch #(  
    // TODO
) (
    input wire clk,
    input wire reset
    // TODO
);

    // TODO

endmodule