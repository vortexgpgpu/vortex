module VX_tex_format #(
    parameter CORE_ID = 0
) (
    // TODO
)   
    // TODO

endmodule