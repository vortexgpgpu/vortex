`include "VX_define.vh"

module VX_tex_mgr (
    input wire clk,
    input wire reset
);

    //--

endmodule
    








