`include "VX_platform.vh"
`include "VX_define.vh"

module VX_tex_pt_addr #(

) (

  );

  // Need to fill in
    
endmodule