// Copyright © 2019-2023
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`include "VX_define.vh"

//Partial product summation result will never exceed 2*N
`define CSA_NO_COUT

module VX_tcu_drl_wallaceTreeMul #(
    parameter N = 8
) (
    input wire [N-1:0] a,
    input wire [N-1:0] b,
    output logic [2*N-1:0] product
);
    wire [2*N-1:0] pp[N-1:0];    //partial products, double width (shifted)
    
    genvar g, h;
    generate
        for(g = 0; g < N; g=g+1) begin: g_pp_loop
            for(h = 0; h < N; h=h+1) begin: g_and_loop
                and a(pp[g][h+g], a[h], b[g]);
            end
            if(g != 0) begin : g_bit_fill
                assign pp[g][g-1:0] = {g{1'b0}};    //fill lower bits with zeros
            end
            assign pp[g][2*N-1:N+g] = {(N-g){1'b0}};    //fill upper bits with zeros 
        end
    endgenerate

    VX_tcu_drl_CSA #(.M(N), .N(2*N)) pp_acc(.Operands(pp), .Sum(product));
endmodule
