`include "VX_rop_define.vh"

// Module for handling memory requests
module VX_rop_mem #(
    // TODO
) (
    input wire clk,
    input wire reset
    // TODO
);

    // TODO

endmodule