`ifndef VORTEX_AFU_VH
`define VORTEX_AFU_VH

`ifndef NOPAE
`include "afu_json_info.vh"
`else
`define PLATFORM_PROVIDES_LOCAL_MEMORY

`ifndef PLATFORM_PARAM_LOCAL_MEMORY_BANKS
`define PLATFORM_PARAM_LOCAL_MEMORY_BANKS 2
`endif

`ifndef PLATFORM_PARAM_LOCAL_MEMORY_ADDR_WIDTH
`define PLATFORM_PARAM_LOCAL_MEMORY_ADDR_WIDTH 26
`endif

`ifndef PLATFORM_PARAM_LOCAL_MEMORY_DATA_WIDTH
`define PLATFORM_PARAM_LOCAL_MEMORY_DATA_WIDTH 512
`endif

`ifndef PLATFORM_PARAM_LOCAL_MEMORY_BURST_CNT_WIDTH
`define PLATFORM_PARAM_LOCAL_MEMORY_BURST_CNT_WIDTH 4
`endif

`define AFU_ACCEL_NAME "vortex_afu"
`define AFU_ACCEL_UUID 128'h35f9452b_25c2_434c_93d5_6f8c60db361c

`define AFU_IMAGE_CMD_MEM_READ 1
`define AFU_IMAGE_CMD_MEM_WRITE 2
`define AFU_IMAGE_CMD_RUN 3
`define AFU_IMAGE_CMD_DCR_WRITE 4
`define AFU_IMAGE_CMD_MAX_VALUE 4

`define AFU_IMAGE_MMIO_CMD_TYPE 10
`define AFU_IMAGE_MMIO_CMD_ARG0 12
`define AFU_IMAGE_MMIO_CMD_ARG1 14
`define AFU_IMAGE_MMIO_CMD_ARG2 16
`define AFU_IMAGE_MMIO_STATUS 18
`define AFU_IMAGE_MMIO_SCOPE_READ 20
`define AFU_IMAGE_MMIO_SCOPE_WRITE 22
`define AFU_IMAGE_MMIO_DEV_CAPS 24
`define AFU_IMAGE_MMIO_ISA_CAPS 26

`define AFU_IMAGE_POWER 0
`define AFU_TOP_IFC "ccip_std_afu_avalon_mm"

`endif // NOPAE

`include "VX_define.vh"
`include "VX_gpu_types.vh"

`endif // VORTEX_AFU_VH
