`include "VX_raster_define.vh"

module VX_raster_rsp_switch #(  
    parameter CORE_ID = 0
    // TODO
) (
    input wire clk,
    input wire reset
    // TODO
);

    // TODO

endmodule