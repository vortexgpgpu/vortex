`ifndef __VORTEX_AFU__
`define __VORTEX_AFU__

`IGNORE_WARNINGS_BEGIN
`include "ccip_if_pkg.sv"
`IGNORE_WARNINGS_END

`define PLATFORM_PROVIDES_LOCAL_MEMORY
`define PLATFORM_PARAM_LOCAL_MEMORY_ADDR_WIDTH      26
`define PLATFORM_PARAM_LOCAL_MEMORY_DATA_WIDTH      512
`define PLATFORM_PARAM_LOCAL_MEMORY_BURST_CNT_WIDTH 4

`IGNORE_WARNINGS_BEGIN
`include "local_mem_cfg_pkg.sv"
`IGNORE_WARNINGS_END

`define AFU_ACCEL_NAME "vortex_afu"
`define AFU_ACCEL_UUID 128'h35f9452b_25c2_434c_93d5_6f8c60db361c

`define AFU_IMAGE_CMD_CSR_READ 4
`define AFU_IMAGE_CMD_CSR_WRITE 5
`define AFU_IMAGE_CMD_MEM_READ 1
`define AFU_IMAGE_CMD_MEM_WRITE 2
`define AFU_IMAGE_CMD_RUN 3
`define AFU_IMAGE_MMIO_CMD_TYPE 10
`define AFU_IMAGE_MMIO_CSR_CORE 24
`define AFU_IMAGE_MMIO_CSR_ADDR 26
`define AFU_IMAGE_MMIO_CSR_DATA 28
`define AFU_IMAGE_MMIO_CSR_READ 30
`define AFU_IMAGE_MMIO_DATA_SIZE 16
`define AFU_IMAGE_MMIO_IO_ADDR 12
`define AFU_IMAGE_MMIO_MEM_ADDR 14
`define AFU_IMAGE_MMIO_SCOPE_READ 20
`define AFU_IMAGE_MMIO_SCOPE_WRITE 22
`define AFU_IMAGE_MMIO_STATUS 18

`define AFU_IMAGE_POWER 0
`define AFU_TOP_IFC "ccip_std_afu_avalon_mm"

`endif