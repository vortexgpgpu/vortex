`include "VX_raster_define.vh"

// Module for triangle setup
//  Description: Perform edge equation computation

module VX_raster_setup #(  
    parameter CORE_ID = 0
    // TODO
) (
    input wire clk,
    input wire reset
    // TODO
);

    // TODO

endmodule