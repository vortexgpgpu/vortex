
`ifndef VX_SCOPE
`define VX_SCOPE

`ifdef SCOPE

`include "scope-defs.vh"

`define SCOPE_ASSIGN(d,s) assign d = s

`else

`define SCOPE_SIGNALS_ISTAGE_TOP_IO
`define SCOPE_SIGNALS_ISTAGE_TOP_BIND
`define SCOPE_SIGNALS_ISTAGE_CLUSTER_IO
`define SCOPE_SIGNALS_ISTAGE_CLUSTER_BIND
`define SCOPE_SIGNALS_ISTAGE_IO
`define SCOPE_SIGNALS_ISTAGE_BIND
`define SCOPE_SIGNALS_ISTAGE_CLUSTER_SELECT(__i__)
`define SCOPE_SIGNALS_ISTAGE_SELECT(__i__)
`define SCOPE_SIGNALS_LSU_TOP_IO
`define SCOPE_SIGNALS_LSU_TOP_BIND
`define SCOPE_SIGNALS_LSU_CLUSTER_IO
`define SCOPE_SIGNALS_LSU_CLUSTER_BIND
`define SCOPE_SIGNALS_LSU_IO
`define SCOPE_SIGNALS_LSU_BIND
`define SCOPE_SIGNALS_LSU_CLUSTER_SELECT(__i__)
`define SCOPE_SIGNALS_LSU_SELECT(__i__)
`define SCOPE_SIGNALS_ISSUE_TOP_IO
`define SCOPE_SIGNALS_ISSUE_TOP_BIND
`define SCOPE_SIGNALS_ISSUE_CLUSTER_IO
`define SCOPE_SIGNALS_ISSUE_CLUSTER_BIND
`define SCOPE_SIGNALS_ISSUE_IO
`define SCOPE_SIGNALS_ISSUE_BIND
`define SCOPE_SIGNALS_ISSUE_CLUSTER_SELECT(__i__)
`define SCOPE_SIGNALS_ISSUE_SELECT(__i__)
`define SCOPE_SIGNALS_EXECUTE_TOP_IO
`define SCOPE_SIGNALS_EXECUTE_TOP_BIND
`define SCOPE_SIGNALS_EXECUTE_CLUSTER_IO
`define SCOPE_SIGNALS_EXECUTE_CLUSTER_BIND
`define SCOPE_SIGNALS_EXECUTE_IO
`define SCOPE_SIGNALS_EXECUTE_BIND
`define SCOPE_SIGNALS_EXECUTE_CLUSTER_SELECT(__i__)
`define SCOPE_SIGNALS_EXECUTE_SELECT(__i__)
`define SCOPE_SIGNALS_BANK_L3_TOP_IO
`define SCOPE_SIGNALS_BANK_L3_TOP_BIND
`define SCOPE_SIGNALS_BANK_L2_TOP_IO
`define SCOPE_SIGNALS_BANK_L2_TOP_BIND
`define SCOPE_SIGNALS_BANK_L1D_TOP_IO
`define SCOPE_SIGNALS_BANK_L1D_TOP_BIND
`define SCOPE_SIGNALS_BANK_L1I_TOP_IO
`define SCOPE_SIGNALS_BANK_L1I_TOP_BIND
`define SCOPE_SIGNALS_BANK_L1S_TOP_IO
`define SCOPE_SIGNALS_BANK_L1S_TOP_BIND
`define SCOPE_SIGNALS_BANK_L2_CLUSTER_IO
`define SCOPE_SIGNALS_BANK_L2_CLUSTER_BIND
`define SCOPE_SIGNALS_BANK_L1D_CLUSTER_IO
`define SCOPE_SIGNALS_BANK_L1D_CLUSTER_BIND
`define SCOPE_SIGNALS_BANK_L1I_CLUSTER_IO
`define SCOPE_SIGNALS_BANK_L1I_CLUSTER_BIND
`define SCOPE_SIGNALS_BANK_L1S_CLUSTER_IO
`define SCOPE_SIGNALS_BANK_L1S_CLUSTER_BIND
`define SCOPE_SIGNALS_BANK_L1D_CORE_IO
`define SCOPE_SIGNALS_BANK_L1D_CORE_BIND
`define SCOPE_SIGNALS_BANK_L1I_CORE_IO
`define SCOPE_SIGNALS_BANK_L1I_CORE_BIND
`define SCOPE_SIGNALS_BANK_L1S_CORE_IO
`define SCOPE_SIGNALS_BANK_L1S_CORE_BIND
`define SCOPE_SIGNALS_BANK_CACHE_IO
`define SCOPE_SIGNALS_BANK_CACHE_BIND
`define SCOPE_SIGNALS_BANK_IO
`define SCOPE_SIGNALS_BANK_BIND
`define SCOPE_SIGNALS_BANK_L2_CLUSTER_SELECT(__i__)
`define SCOPE_SIGNALS_BANK_L1D_CLUSTER_SELECT(__i__)
`define SCOPE_SIGNALS_BANK_L1I_CLUSTER_SELECT(__i__)
`define SCOPE_SIGNALS_BANK_L1S_CLUSTER_SELECT(__i__)
`define SCOPE_SIGNALS_BANK_L1D_CORE_SELECT(__i__)
`define SCOPE_SIGNALS_BANK_L1I_CORE_SELECT(__i__)
`define SCOPE_SIGNALS_BANK_L1S_CORE_SELECT(__i__)
`define SCOPE_SIGNALS_BANK_L3_CACHE_BIND
`define SCOPE_SIGNALS_BANK_L2_CACHE_BIND
`define SCOPE_SIGNALS_BANK_L1D_CACHE_BIND
`define SCOPE_SIGNALS_BANK_L1I_CACHE_BIND
`define SCOPE_SIGNALS_BANK_L1S_CACHE_BIND
`define SCOPE_SIGNALS_BANK_SELECT(__i__)
`define SCOPE_ASSIGN(d,s)

`endif
`endif