`ifndef VX_CACHE_TYPES_VH
`define VX_CACHE_TYPES_VH

`include "VX_cache_define.vh"

package VX_cache_types;

`define _ICACHE_TAG_WIDTH       (`ICACHE_NOSM_TAG_WIDTH + `ARB_SEL_BITS(`NUM_CORES, `UP(`NUM_ICACHES)))
`ifdef ICACHE_ENABLE
`define _ICACHE_MEM_TAG_WIDTH   `CACHE_MEM_TAG_WIDTH(`ICACHE_MSHR_SIZE, `ICACHE_NUM_BANKS)
`else
`define _ICACHE_MEM_TAG_WIDTH   `CACHE_BYPASS_TAG_WIDTH(`ICACHE_NUM_REQS, `ICACHE_LINE_SIZE, `ICACHE_WORD_SIZE, `_ICACHE_TAG_WIDTH)
`endif
localparam ICACHE_MEM_TAG_WIDTH = (`_ICACHE_MEM_TAG_WIDTH + `ARB_SEL_BITS(`UP(`NUM_ICACHES), 1));

`define DCACHE_NOSM_TAG_WIDTH   (`DCACHE_TAG_WIDTH - `SM_ENABLED)
`define _DCACHE_NOSM_TAG_WIDTH  (`DCACHE_NOSM_TAG_WIDTH + `ARB_SEL_BITS(`NUM_CORES, `UP(`NUM_DCACHES)))
`ifdef DCACHE_ENABLE
`define _DCACHE_MEM_TAG_WIDTH   `CACHE_NC_MEM_TAG_WIDTH(`DCACHE_MSHR_SIZE, `DCACHE_NUM_BANKS, `DCACHE_NUM_REQS, `DCACHE_LINE_SIZE, `DCACHE_WORD_SIZE, `_DCACHE_NOSM_TAG_WIDTH)
`else
`define _DCACHE_MEM_TAG_WIDTH   `CACHE_NC_BYPASS_TAG_WIDTH(`DCACHE_NUM_REQS, `DCACHE_LINE_SIZE, `DCACHE_WORD_SIZE, `DCACHE_TAG_WIDTH)
`endif
localparam DCACHE_MEM_TAG_WIDTH = (`_DCACHE_MEM_TAG_WIDTH + `ARB_SEL_BITS(`UP(`NUM_DCACHES), 1));

`ifdef L2_ENABLE
`define _L2_MEM_TAG_WIDTH       `CACHE_NC_MEM_TAG_WIDTH(`L2_MSHR_SIZE, `L2_NUM_BANKS, `L2_NUM_REQS, `L2_LINE_SIZE, `L2_WORD_SIZE, `L2_TAG_WIDTH)
`else
`define _L2_MEM_TAG_WIDTH       `CACHE_NC_BYPASS_TAG_WIDTH(`L2_NUM_REQS, `L2_LINE_SIZE, `L2_WORD_SIZE, `L2_TAG_WIDTH)
`endif
localparam L2_MEM_TAG_WIDTH = `_L2_MEM_TAG_WIDTH;

`ifdef L3_ENABLE
`define _L3_MEM_TAG_WIDTH       `CACHE_NC_MEM_TAG_WIDTH(`L3_MSHR_SIZE, `L3_NUM_BANKS, `L3_NUM_REQS, `L3_LINE_SIZE, `L3_WORD_SIZE, `L3_TAG_WIDTH)
`else
`define _L3_MEM_TAG_WIDTH       `CACHE_NC_BYPASS_TAG_WIDTH(`L3_NUM_REQS, `L3_LINE_SIZE, `L3_WORD_SIZE, `L3_TAG_WIDTH)
`endif
localparam L3_MEM_TAG_WIDTH = `_L3_MEM_TAG_WIDTH;

endpackage

`endif
