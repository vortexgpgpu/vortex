`ifndef VX_RASTER_DEFINE_VH
`define VX_RASTER_DEFINE_VH

`include "VX_define.vh"
`include "VX_raster_types.vh"

`IGNORE_WARNINGS_BEGIN
import VX_raster_types::*;
`IGNORE_WARNINGS_END

`endif
