`include "VX_raster_define.vh"

// Module for primitive fetch
//  Descrption: Performs strided fetch
//  of primitive data from the buffer

module VX_raster_fetch #(  
    parameter CORE_ID = 0
    // TODO
) (
    input wire clk,
    input wire reset
    // TODO
);

    // TODO
    `UNUSED_VAR (clk)
    `UNUSED_VAR (reset)

endmodule